`ifndef __EPU_def__
`define __EPU_def__

    `define EPU_DATA_BITS 32
    `define EPU_ADDR_BITS 17

`endif