`ifndef __CACHEFL__
`define __CACHEFL__

module cachefilter (
    input  [31:0] addr_i,
    output        volatile_o
);

    // assign volatile_o = ()

endmodule
`endif