# 
#              Synchronous High Speed Single Port SRAM Compiler 
# 
#                    UMC 0.18um GenericII Logic Process
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : SUMA180_384X32X1BM4
#       Words            : 384
#       Bits             : 32
#       Byte-Write       : 1
#       Aspect Ratio     : 4
#       Output Loading   : 0.5  (pf)
#       Data Slew        : 0.5  (ns)
#       CK Slew          : 0.5  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2022/01/11 11:39:30
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO SUMA180_384X32X1BM4
CLASS BLOCK ;
FOREIGN SUMA180_384X32X1BM4 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 1899.060 BY 166.880 ;
SYMMETRY x y r90 ;
SITE core ;
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 1897.940 129.700 1899.060 132.940 ;
  LAYER metal3 ;
  RECT 1897.940 129.700 1899.060 132.940 ;
  LAYER metal2 ;
  RECT 1897.940 129.700 1899.060 132.940 ;
  LAYER metal1 ;
  RECT 1897.940 129.700 1899.060 132.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1897.940 121.860 1899.060 125.100 ;
  LAYER metal3 ;
  RECT 1897.940 121.860 1899.060 125.100 ;
  LAYER metal2 ;
  RECT 1897.940 121.860 1899.060 125.100 ;
  LAYER metal1 ;
  RECT 1897.940 121.860 1899.060 125.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1897.940 114.020 1899.060 117.260 ;
  LAYER metal3 ;
  RECT 1897.940 114.020 1899.060 117.260 ;
  LAYER metal2 ;
  RECT 1897.940 114.020 1899.060 117.260 ;
  LAYER metal1 ;
  RECT 1897.940 114.020 1899.060 117.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1897.940 106.180 1899.060 109.420 ;
  LAYER metal3 ;
  RECT 1897.940 106.180 1899.060 109.420 ;
  LAYER metal2 ;
  RECT 1897.940 106.180 1899.060 109.420 ;
  LAYER metal1 ;
  RECT 1897.940 106.180 1899.060 109.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1897.940 98.340 1899.060 101.580 ;
  LAYER metal3 ;
  RECT 1897.940 98.340 1899.060 101.580 ;
  LAYER metal2 ;
  RECT 1897.940 98.340 1899.060 101.580 ;
  LAYER metal1 ;
  RECT 1897.940 98.340 1899.060 101.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1897.940 90.500 1899.060 93.740 ;
  LAYER metal3 ;
  RECT 1897.940 90.500 1899.060 93.740 ;
  LAYER metal2 ;
  RECT 1897.940 90.500 1899.060 93.740 ;
  LAYER metal1 ;
  RECT 1897.940 90.500 1899.060 93.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1897.940 51.300 1899.060 54.540 ;
  LAYER metal3 ;
  RECT 1897.940 51.300 1899.060 54.540 ;
  LAYER metal2 ;
  RECT 1897.940 51.300 1899.060 54.540 ;
  LAYER metal1 ;
  RECT 1897.940 51.300 1899.060 54.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1897.940 43.460 1899.060 46.700 ;
  LAYER metal3 ;
  RECT 1897.940 43.460 1899.060 46.700 ;
  LAYER metal2 ;
  RECT 1897.940 43.460 1899.060 46.700 ;
  LAYER metal1 ;
  RECT 1897.940 43.460 1899.060 46.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1897.940 35.620 1899.060 38.860 ;
  LAYER metal3 ;
  RECT 1897.940 35.620 1899.060 38.860 ;
  LAYER metal2 ;
  RECT 1897.940 35.620 1899.060 38.860 ;
  LAYER metal1 ;
  RECT 1897.940 35.620 1899.060 38.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1897.940 27.780 1899.060 31.020 ;
  LAYER metal3 ;
  RECT 1897.940 27.780 1899.060 31.020 ;
  LAYER metal2 ;
  RECT 1897.940 27.780 1899.060 31.020 ;
  LAYER metal1 ;
  RECT 1897.940 27.780 1899.060 31.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1897.940 19.940 1899.060 23.180 ;
  LAYER metal3 ;
  RECT 1897.940 19.940 1899.060 23.180 ;
  LAYER metal2 ;
  RECT 1897.940 19.940 1899.060 23.180 ;
  LAYER metal1 ;
  RECT 1897.940 19.940 1899.060 23.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1897.940 12.100 1899.060 15.340 ;
  LAYER metal3 ;
  RECT 1897.940 12.100 1899.060 15.340 ;
  LAYER metal2 ;
  RECT 1897.940 12.100 1899.060 15.340 ;
  LAYER metal1 ;
  RECT 1897.940 12.100 1899.060 15.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal3 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal2 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal1 ;
  RECT 0.000 129.700 1.120 132.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal3 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal2 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal1 ;
  RECT 0.000 121.860 1.120 125.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal3 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal2 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal1 ;
  RECT 0.000 114.020 1.120 117.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal3 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal2 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal1 ;
  RECT 0.000 106.180 1.120 109.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal3 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal2 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal1 ;
  RECT 0.000 98.340 1.120 101.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal3 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal2 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal1 ;
  RECT 0.000 90.500 1.120 93.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal3 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal2 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal1 ;
  RECT 0.000 51.300 1.120 54.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal3 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal2 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal1 ;
  RECT 0.000 43.460 1.120 46.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal3 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal2 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal1 ;
  RECT 0.000 35.620 1.120 38.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal3 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal2 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal1 ;
  RECT 0.000 27.780 1.120 31.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal3 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal2 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal1 ;
  RECT 0.000 19.940 1.120 23.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal3 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal2 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal1 ;
  RECT 0.000 12.100 1.120 15.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1878.380 165.760 1881.920 166.880 ;
  LAYER metal3 ;
  RECT 1878.380 165.760 1881.920 166.880 ;
  LAYER metal2 ;
  RECT 1878.380 165.760 1881.920 166.880 ;
  LAYER metal1 ;
  RECT 1878.380 165.760 1881.920 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1869.700 165.760 1873.240 166.880 ;
  LAYER metal3 ;
  RECT 1869.700 165.760 1873.240 166.880 ;
  LAYER metal2 ;
  RECT 1869.700 165.760 1873.240 166.880 ;
  LAYER metal1 ;
  RECT 1869.700 165.760 1873.240 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1861.020 165.760 1864.560 166.880 ;
  LAYER metal3 ;
  RECT 1861.020 165.760 1864.560 166.880 ;
  LAYER metal2 ;
  RECT 1861.020 165.760 1864.560 166.880 ;
  LAYER metal1 ;
  RECT 1861.020 165.760 1864.560 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1852.340 165.760 1855.880 166.880 ;
  LAYER metal3 ;
  RECT 1852.340 165.760 1855.880 166.880 ;
  LAYER metal2 ;
  RECT 1852.340 165.760 1855.880 166.880 ;
  LAYER metal1 ;
  RECT 1852.340 165.760 1855.880 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1843.660 165.760 1847.200 166.880 ;
  LAYER metal3 ;
  RECT 1843.660 165.760 1847.200 166.880 ;
  LAYER metal2 ;
  RECT 1843.660 165.760 1847.200 166.880 ;
  LAYER metal1 ;
  RECT 1843.660 165.760 1847.200 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1834.980 165.760 1838.520 166.880 ;
  LAYER metal3 ;
  RECT 1834.980 165.760 1838.520 166.880 ;
  LAYER metal2 ;
  RECT 1834.980 165.760 1838.520 166.880 ;
  LAYER metal1 ;
  RECT 1834.980 165.760 1838.520 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1791.580 165.760 1795.120 166.880 ;
  LAYER metal3 ;
  RECT 1791.580 165.760 1795.120 166.880 ;
  LAYER metal2 ;
  RECT 1791.580 165.760 1795.120 166.880 ;
  LAYER metal1 ;
  RECT 1791.580 165.760 1795.120 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1782.900 165.760 1786.440 166.880 ;
  LAYER metal3 ;
  RECT 1782.900 165.760 1786.440 166.880 ;
  LAYER metal2 ;
  RECT 1782.900 165.760 1786.440 166.880 ;
  LAYER metal1 ;
  RECT 1782.900 165.760 1786.440 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1774.220 165.760 1777.760 166.880 ;
  LAYER metal3 ;
  RECT 1774.220 165.760 1777.760 166.880 ;
  LAYER metal2 ;
  RECT 1774.220 165.760 1777.760 166.880 ;
  LAYER metal1 ;
  RECT 1774.220 165.760 1777.760 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1765.540 165.760 1769.080 166.880 ;
  LAYER metal3 ;
  RECT 1765.540 165.760 1769.080 166.880 ;
  LAYER metal2 ;
  RECT 1765.540 165.760 1769.080 166.880 ;
  LAYER metal1 ;
  RECT 1765.540 165.760 1769.080 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1756.860 165.760 1760.400 166.880 ;
  LAYER metal3 ;
  RECT 1756.860 165.760 1760.400 166.880 ;
  LAYER metal2 ;
  RECT 1756.860 165.760 1760.400 166.880 ;
  LAYER metal1 ;
  RECT 1756.860 165.760 1760.400 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1748.180 165.760 1751.720 166.880 ;
  LAYER metal3 ;
  RECT 1748.180 165.760 1751.720 166.880 ;
  LAYER metal2 ;
  RECT 1748.180 165.760 1751.720 166.880 ;
  LAYER metal1 ;
  RECT 1748.180 165.760 1751.720 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1704.780 165.760 1708.320 166.880 ;
  LAYER metal3 ;
  RECT 1704.780 165.760 1708.320 166.880 ;
  LAYER metal2 ;
  RECT 1704.780 165.760 1708.320 166.880 ;
  LAYER metal1 ;
  RECT 1704.780 165.760 1708.320 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1696.100 165.760 1699.640 166.880 ;
  LAYER metal3 ;
  RECT 1696.100 165.760 1699.640 166.880 ;
  LAYER metal2 ;
  RECT 1696.100 165.760 1699.640 166.880 ;
  LAYER metal1 ;
  RECT 1696.100 165.760 1699.640 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1687.420 165.760 1690.960 166.880 ;
  LAYER metal3 ;
  RECT 1687.420 165.760 1690.960 166.880 ;
  LAYER metal2 ;
  RECT 1687.420 165.760 1690.960 166.880 ;
  LAYER metal1 ;
  RECT 1687.420 165.760 1690.960 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1678.740 165.760 1682.280 166.880 ;
  LAYER metal3 ;
  RECT 1678.740 165.760 1682.280 166.880 ;
  LAYER metal2 ;
  RECT 1678.740 165.760 1682.280 166.880 ;
  LAYER metal1 ;
  RECT 1678.740 165.760 1682.280 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1670.060 165.760 1673.600 166.880 ;
  LAYER metal3 ;
  RECT 1670.060 165.760 1673.600 166.880 ;
  LAYER metal2 ;
  RECT 1670.060 165.760 1673.600 166.880 ;
  LAYER metal1 ;
  RECT 1670.060 165.760 1673.600 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1661.380 165.760 1664.920 166.880 ;
  LAYER metal3 ;
  RECT 1661.380 165.760 1664.920 166.880 ;
  LAYER metal2 ;
  RECT 1661.380 165.760 1664.920 166.880 ;
  LAYER metal1 ;
  RECT 1661.380 165.760 1664.920 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1617.980 165.760 1621.520 166.880 ;
  LAYER metal3 ;
  RECT 1617.980 165.760 1621.520 166.880 ;
  LAYER metal2 ;
  RECT 1617.980 165.760 1621.520 166.880 ;
  LAYER metal1 ;
  RECT 1617.980 165.760 1621.520 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1609.300 165.760 1612.840 166.880 ;
  LAYER metal3 ;
  RECT 1609.300 165.760 1612.840 166.880 ;
  LAYER metal2 ;
  RECT 1609.300 165.760 1612.840 166.880 ;
  LAYER metal1 ;
  RECT 1609.300 165.760 1612.840 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1600.620 165.760 1604.160 166.880 ;
  LAYER metal3 ;
  RECT 1600.620 165.760 1604.160 166.880 ;
  LAYER metal2 ;
  RECT 1600.620 165.760 1604.160 166.880 ;
  LAYER metal1 ;
  RECT 1600.620 165.760 1604.160 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1591.940 165.760 1595.480 166.880 ;
  LAYER metal3 ;
  RECT 1591.940 165.760 1595.480 166.880 ;
  LAYER metal2 ;
  RECT 1591.940 165.760 1595.480 166.880 ;
  LAYER metal1 ;
  RECT 1591.940 165.760 1595.480 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1583.260 165.760 1586.800 166.880 ;
  LAYER metal3 ;
  RECT 1583.260 165.760 1586.800 166.880 ;
  LAYER metal2 ;
  RECT 1583.260 165.760 1586.800 166.880 ;
  LAYER metal1 ;
  RECT 1583.260 165.760 1586.800 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1574.580 165.760 1578.120 166.880 ;
  LAYER metal3 ;
  RECT 1574.580 165.760 1578.120 166.880 ;
  LAYER metal2 ;
  RECT 1574.580 165.760 1578.120 166.880 ;
  LAYER metal1 ;
  RECT 1574.580 165.760 1578.120 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1531.180 165.760 1534.720 166.880 ;
  LAYER metal3 ;
  RECT 1531.180 165.760 1534.720 166.880 ;
  LAYER metal2 ;
  RECT 1531.180 165.760 1534.720 166.880 ;
  LAYER metal1 ;
  RECT 1531.180 165.760 1534.720 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1522.500 165.760 1526.040 166.880 ;
  LAYER metal3 ;
  RECT 1522.500 165.760 1526.040 166.880 ;
  LAYER metal2 ;
  RECT 1522.500 165.760 1526.040 166.880 ;
  LAYER metal1 ;
  RECT 1522.500 165.760 1526.040 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1513.820 165.760 1517.360 166.880 ;
  LAYER metal3 ;
  RECT 1513.820 165.760 1517.360 166.880 ;
  LAYER metal2 ;
  RECT 1513.820 165.760 1517.360 166.880 ;
  LAYER metal1 ;
  RECT 1513.820 165.760 1517.360 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1505.140 165.760 1508.680 166.880 ;
  LAYER metal3 ;
  RECT 1505.140 165.760 1508.680 166.880 ;
  LAYER metal2 ;
  RECT 1505.140 165.760 1508.680 166.880 ;
  LAYER metal1 ;
  RECT 1505.140 165.760 1508.680 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1496.460 165.760 1500.000 166.880 ;
  LAYER metal3 ;
  RECT 1496.460 165.760 1500.000 166.880 ;
  LAYER metal2 ;
  RECT 1496.460 165.760 1500.000 166.880 ;
  LAYER metal1 ;
  RECT 1496.460 165.760 1500.000 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1487.780 165.760 1491.320 166.880 ;
  LAYER metal3 ;
  RECT 1487.780 165.760 1491.320 166.880 ;
  LAYER metal2 ;
  RECT 1487.780 165.760 1491.320 166.880 ;
  LAYER metal1 ;
  RECT 1487.780 165.760 1491.320 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1444.380 165.760 1447.920 166.880 ;
  LAYER metal3 ;
  RECT 1444.380 165.760 1447.920 166.880 ;
  LAYER metal2 ;
  RECT 1444.380 165.760 1447.920 166.880 ;
  LAYER metal1 ;
  RECT 1444.380 165.760 1447.920 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1435.700 165.760 1439.240 166.880 ;
  LAYER metal3 ;
  RECT 1435.700 165.760 1439.240 166.880 ;
  LAYER metal2 ;
  RECT 1435.700 165.760 1439.240 166.880 ;
  LAYER metal1 ;
  RECT 1435.700 165.760 1439.240 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1427.020 165.760 1430.560 166.880 ;
  LAYER metal3 ;
  RECT 1427.020 165.760 1430.560 166.880 ;
  LAYER metal2 ;
  RECT 1427.020 165.760 1430.560 166.880 ;
  LAYER metal1 ;
  RECT 1427.020 165.760 1430.560 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1418.340 165.760 1421.880 166.880 ;
  LAYER metal3 ;
  RECT 1418.340 165.760 1421.880 166.880 ;
  LAYER metal2 ;
  RECT 1418.340 165.760 1421.880 166.880 ;
  LAYER metal1 ;
  RECT 1418.340 165.760 1421.880 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1409.660 165.760 1413.200 166.880 ;
  LAYER metal3 ;
  RECT 1409.660 165.760 1413.200 166.880 ;
  LAYER metal2 ;
  RECT 1409.660 165.760 1413.200 166.880 ;
  LAYER metal1 ;
  RECT 1409.660 165.760 1413.200 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1400.980 165.760 1404.520 166.880 ;
  LAYER metal3 ;
  RECT 1400.980 165.760 1404.520 166.880 ;
  LAYER metal2 ;
  RECT 1400.980 165.760 1404.520 166.880 ;
  LAYER metal1 ;
  RECT 1400.980 165.760 1404.520 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1357.580 165.760 1361.120 166.880 ;
  LAYER metal3 ;
  RECT 1357.580 165.760 1361.120 166.880 ;
  LAYER metal2 ;
  RECT 1357.580 165.760 1361.120 166.880 ;
  LAYER metal1 ;
  RECT 1357.580 165.760 1361.120 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1348.900 165.760 1352.440 166.880 ;
  LAYER metal3 ;
  RECT 1348.900 165.760 1352.440 166.880 ;
  LAYER metal2 ;
  RECT 1348.900 165.760 1352.440 166.880 ;
  LAYER metal1 ;
  RECT 1348.900 165.760 1352.440 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1340.220 165.760 1343.760 166.880 ;
  LAYER metal3 ;
  RECT 1340.220 165.760 1343.760 166.880 ;
  LAYER metal2 ;
  RECT 1340.220 165.760 1343.760 166.880 ;
  LAYER metal1 ;
  RECT 1340.220 165.760 1343.760 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1331.540 165.760 1335.080 166.880 ;
  LAYER metal3 ;
  RECT 1331.540 165.760 1335.080 166.880 ;
  LAYER metal2 ;
  RECT 1331.540 165.760 1335.080 166.880 ;
  LAYER metal1 ;
  RECT 1331.540 165.760 1335.080 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1322.860 165.760 1326.400 166.880 ;
  LAYER metal3 ;
  RECT 1322.860 165.760 1326.400 166.880 ;
  LAYER metal2 ;
  RECT 1322.860 165.760 1326.400 166.880 ;
  LAYER metal1 ;
  RECT 1322.860 165.760 1326.400 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1314.180 165.760 1317.720 166.880 ;
  LAYER metal3 ;
  RECT 1314.180 165.760 1317.720 166.880 ;
  LAYER metal2 ;
  RECT 1314.180 165.760 1317.720 166.880 ;
  LAYER metal1 ;
  RECT 1314.180 165.760 1317.720 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1270.780 165.760 1274.320 166.880 ;
  LAYER metal3 ;
  RECT 1270.780 165.760 1274.320 166.880 ;
  LAYER metal2 ;
  RECT 1270.780 165.760 1274.320 166.880 ;
  LAYER metal1 ;
  RECT 1270.780 165.760 1274.320 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1262.100 165.760 1265.640 166.880 ;
  LAYER metal3 ;
  RECT 1262.100 165.760 1265.640 166.880 ;
  LAYER metal2 ;
  RECT 1262.100 165.760 1265.640 166.880 ;
  LAYER metal1 ;
  RECT 1262.100 165.760 1265.640 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1253.420 165.760 1256.960 166.880 ;
  LAYER metal3 ;
  RECT 1253.420 165.760 1256.960 166.880 ;
  LAYER metal2 ;
  RECT 1253.420 165.760 1256.960 166.880 ;
  LAYER metal1 ;
  RECT 1253.420 165.760 1256.960 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1244.740 165.760 1248.280 166.880 ;
  LAYER metal3 ;
  RECT 1244.740 165.760 1248.280 166.880 ;
  LAYER metal2 ;
  RECT 1244.740 165.760 1248.280 166.880 ;
  LAYER metal1 ;
  RECT 1244.740 165.760 1248.280 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1236.060 165.760 1239.600 166.880 ;
  LAYER metal3 ;
  RECT 1236.060 165.760 1239.600 166.880 ;
  LAYER metal2 ;
  RECT 1236.060 165.760 1239.600 166.880 ;
  LAYER metal1 ;
  RECT 1236.060 165.760 1239.600 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1227.380 165.760 1230.920 166.880 ;
  LAYER metal3 ;
  RECT 1227.380 165.760 1230.920 166.880 ;
  LAYER metal2 ;
  RECT 1227.380 165.760 1230.920 166.880 ;
  LAYER metal1 ;
  RECT 1227.380 165.760 1230.920 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1183.980 165.760 1187.520 166.880 ;
  LAYER metal3 ;
  RECT 1183.980 165.760 1187.520 166.880 ;
  LAYER metal2 ;
  RECT 1183.980 165.760 1187.520 166.880 ;
  LAYER metal1 ;
  RECT 1183.980 165.760 1187.520 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1175.300 165.760 1178.840 166.880 ;
  LAYER metal3 ;
  RECT 1175.300 165.760 1178.840 166.880 ;
  LAYER metal2 ;
  RECT 1175.300 165.760 1178.840 166.880 ;
  LAYER metal1 ;
  RECT 1175.300 165.760 1178.840 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1166.620 165.760 1170.160 166.880 ;
  LAYER metal3 ;
  RECT 1166.620 165.760 1170.160 166.880 ;
  LAYER metal2 ;
  RECT 1166.620 165.760 1170.160 166.880 ;
  LAYER metal1 ;
  RECT 1166.620 165.760 1170.160 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1157.940 165.760 1161.480 166.880 ;
  LAYER metal3 ;
  RECT 1157.940 165.760 1161.480 166.880 ;
  LAYER metal2 ;
  RECT 1157.940 165.760 1161.480 166.880 ;
  LAYER metal1 ;
  RECT 1157.940 165.760 1161.480 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1149.260 165.760 1152.800 166.880 ;
  LAYER metal3 ;
  RECT 1149.260 165.760 1152.800 166.880 ;
  LAYER metal2 ;
  RECT 1149.260 165.760 1152.800 166.880 ;
  LAYER metal1 ;
  RECT 1149.260 165.760 1152.800 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1140.580 165.760 1144.120 166.880 ;
  LAYER metal3 ;
  RECT 1140.580 165.760 1144.120 166.880 ;
  LAYER metal2 ;
  RECT 1140.580 165.760 1144.120 166.880 ;
  LAYER metal1 ;
  RECT 1140.580 165.760 1144.120 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1097.180 165.760 1100.720 166.880 ;
  LAYER metal3 ;
  RECT 1097.180 165.760 1100.720 166.880 ;
  LAYER metal2 ;
  RECT 1097.180 165.760 1100.720 166.880 ;
  LAYER metal1 ;
  RECT 1097.180 165.760 1100.720 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1088.500 165.760 1092.040 166.880 ;
  LAYER metal3 ;
  RECT 1088.500 165.760 1092.040 166.880 ;
  LAYER metal2 ;
  RECT 1088.500 165.760 1092.040 166.880 ;
  LAYER metal1 ;
  RECT 1088.500 165.760 1092.040 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1079.820 165.760 1083.360 166.880 ;
  LAYER metal3 ;
  RECT 1079.820 165.760 1083.360 166.880 ;
  LAYER metal2 ;
  RECT 1079.820 165.760 1083.360 166.880 ;
  LAYER metal1 ;
  RECT 1079.820 165.760 1083.360 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1071.140 165.760 1074.680 166.880 ;
  LAYER metal3 ;
  RECT 1071.140 165.760 1074.680 166.880 ;
  LAYER metal2 ;
  RECT 1071.140 165.760 1074.680 166.880 ;
  LAYER metal1 ;
  RECT 1071.140 165.760 1074.680 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1062.460 165.760 1066.000 166.880 ;
  LAYER metal3 ;
  RECT 1062.460 165.760 1066.000 166.880 ;
  LAYER metal2 ;
  RECT 1062.460 165.760 1066.000 166.880 ;
  LAYER metal1 ;
  RECT 1062.460 165.760 1066.000 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1053.780 165.760 1057.320 166.880 ;
  LAYER metal3 ;
  RECT 1053.780 165.760 1057.320 166.880 ;
  LAYER metal2 ;
  RECT 1053.780 165.760 1057.320 166.880 ;
  LAYER metal1 ;
  RECT 1053.780 165.760 1057.320 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1010.380 165.760 1013.920 166.880 ;
  LAYER metal3 ;
  RECT 1010.380 165.760 1013.920 166.880 ;
  LAYER metal2 ;
  RECT 1010.380 165.760 1013.920 166.880 ;
  LAYER metal1 ;
  RECT 1010.380 165.760 1013.920 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1001.700 165.760 1005.240 166.880 ;
  LAYER metal3 ;
  RECT 1001.700 165.760 1005.240 166.880 ;
  LAYER metal2 ;
  RECT 1001.700 165.760 1005.240 166.880 ;
  LAYER metal1 ;
  RECT 1001.700 165.760 1005.240 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 993.020 165.760 996.560 166.880 ;
  LAYER metal3 ;
  RECT 993.020 165.760 996.560 166.880 ;
  LAYER metal2 ;
  RECT 993.020 165.760 996.560 166.880 ;
  LAYER metal1 ;
  RECT 993.020 165.760 996.560 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 984.340 165.760 987.880 166.880 ;
  LAYER metal3 ;
  RECT 984.340 165.760 987.880 166.880 ;
  LAYER metal2 ;
  RECT 984.340 165.760 987.880 166.880 ;
  LAYER metal1 ;
  RECT 984.340 165.760 987.880 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 975.660 165.760 979.200 166.880 ;
  LAYER metal3 ;
  RECT 975.660 165.760 979.200 166.880 ;
  LAYER metal2 ;
  RECT 975.660 165.760 979.200 166.880 ;
  LAYER metal1 ;
  RECT 975.660 165.760 979.200 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 966.980 165.760 970.520 166.880 ;
  LAYER metal3 ;
  RECT 966.980 165.760 970.520 166.880 ;
  LAYER metal2 ;
  RECT 966.980 165.760 970.520 166.880 ;
  LAYER metal1 ;
  RECT 966.980 165.760 970.520 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 923.580 165.760 927.120 166.880 ;
  LAYER metal3 ;
  RECT 923.580 165.760 927.120 166.880 ;
  LAYER metal2 ;
  RECT 923.580 165.760 927.120 166.880 ;
  LAYER metal1 ;
  RECT 923.580 165.760 927.120 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 914.900 165.760 918.440 166.880 ;
  LAYER metal3 ;
  RECT 914.900 165.760 918.440 166.880 ;
  LAYER metal2 ;
  RECT 914.900 165.760 918.440 166.880 ;
  LAYER metal1 ;
  RECT 914.900 165.760 918.440 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 906.220 165.760 909.760 166.880 ;
  LAYER metal3 ;
  RECT 906.220 165.760 909.760 166.880 ;
  LAYER metal2 ;
  RECT 906.220 165.760 909.760 166.880 ;
  LAYER metal1 ;
  RECT 906.220 165.760 909.760 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 897.540 165.760 901.080 166.880 ;
  LAYER metal3 ;
  RECT 897.540 165.760 901.080 166.880 ;
  LAYER metal2 ;
  RECT 897.540 165.760 901.080 166.880 ;
  LAYER metal1 ;
  RECT 897.540 165.760 901.080 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 888.860 165.760 892.400 166.880 ;
  LAYER metal3 ;
  RECT 888.860 165.760 892.400 166.880 ;
  LAYER metal2 ;
  RECT 888.860 165.760 892.400 166.880 ;
  LAYER metal1 ;
  RECT 888.860 165.760 892.400 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 880.180 165.760 883.720 166.880 ;
  LAYER metal3 ;
  RECT 880.180 165.760 883.720 166.880 ;
  LAYER metal2 ;
  RECT 880.180 165.760 883.720 166.880 ;
  LAYER metal1 ;
  RECT 880.180 165.760 883.720 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 836.780 165.760 840.320 166.880 ;
  LAYER metal3 ;
  RECT 836.780 165.760 840.320 166.880 ;
  LAYER metal2 ;
  RECT 836.780 165.760 840.320 166.880 ;
  LAYER metal1 ;
  RECT 836.780 165.760 840.320 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 828.100 165.760 831.640 166.880 ;
  LAYER metal3 ;
  RECT 828.100 165.760 831.640 166.880 ;
  LAYER metal2 ;
  RECT 828.100 165.760 831.640 166.880 ;
  LAYER metal1 ;
  RECT 828.100 165.760 831.640 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 819.420 165.760 822.960 166.880 ;
  LAYER metal3 ;
  RECT 819.420 165.760 822.960 166.880 ;
  LAYER metal2 ;
  RECT 819.420 165.760 822.960 166.880 ;
  LAYER metal1 ;
  RECT 819.420 165.760 822.960 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 810.740 165.760 814.280 166.880 ;
  LAYER metal3 ;
  RECT 810.740 165.760 814.280 166.880 ;
  LAYER metal2 ;
  RECT 810.740 165.760 814.280 166.880 ;
  LAYER metal1 ;
  RECT 810.740 165.760 814.280 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 802.060 165.760 805.600 166.880 ;
  LAYER metal3 ;
  RECT 802.060 165.760 805.600 166.880 ;
  LAYER metal2 ;
  RECT 802.060 165.760 805.600 166.880 ;
  LAYER metal1 ;
  RECT 802.060 165.760 805.600 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 793.380 165.760 796.920 166.880 ;
  LAYER metal3 ;
  RECT 793.380 165.760 796.920 166.880 ;
  LAYER metal2 ;
  RECT 793.380 165.760 796.920 166.880 ;
  LAYER metal1 ;
  RECT 793.380 165.760 796.920 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 749.980 165.760 753.520 166.880 ;
  LAYER metal3 ;
  RECT 749.980 165.760 753.520 166.880 ;
  LAYER metal2 ;
  RECT 749.980 165.760 753.520 166.880 ;
  LAYER metal1 ;
  RECT 749.980 165.760 753.520 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 741.300 165.760 744.840 166.880 ;
  LAYER metal3 ;
  RECT 741.300 165.760 744.840 166.880 ;
  LAYER metal2 ;
  RECT 741.300 165.760 744.840 166.880 ;
  LAYER metal1 ;
  RECT 741.300 165.760 744.840 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 732.620 165.760 736.160 166.880 ;
  LAYER metal3 ;
  RECT 732.620 165.760 736.160 166.880 ;
  LAYER metal2 ;
  RECT 732.620 165.760 736.160 166.880 ;
  LAYER metal1 ;
  RECT 732.620 165.760 736.160 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 723.940 165.760 727.480 166.880 ;
  LAYER metal3 ;
  RECT 723.940 165.760 727.480 166.880 ;
  LAYER metal2 ;
  RECT 723.940 165.760 727.480 166.880 ;
  LAYER metal1 ;
  RECT 723.940 165.760 727.480 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 715.260 165.760 718.800 166.880 ;
  LAYER metal3 ;
  RECT 715.260 165.760 718.800 166.880 ;
  LAYER metal2 ;
  RECT 715.260 165.760 718.800 166.880 ;
  LAYER metal1 ;
  RECT 715.260 165.760 718.800 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 706.580 165.760 710.120 166.880 ;
  LAYER metal3 ;
  RECT 706.580 165.760 710.120 166.880 ;
  LAYER metal2 ;
  RECT 706.580 165.760 710.120 166.880 ;
  LAYER metal1 ;
  RECT 706.580 165.760 710.120 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 663.180 165.760 666.720 166.880 ;
  LAYER metal3 ;
  RECT 663.180 165.760 666.720 166.880 ;
  LAYER metal2 ;
  RECT 663.180 165.760 666.720 166.880 ;
  LAYER metal1 ;
  RECT 663.180 165.760 666.720 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 654.500 165.760 658.040 166.880 ;
  LAYER metal3 ;
  RECT 654.500 165.760 658.040 166.880 ;
  LAYER metal2 ;
  RECT 654.500 165.760 658.040 166.880 ;
  LAYER metal1 ;
  RECT 654.500 165.760 658.040 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 645.820 165.760 649.360 166.880 ;
  LAYER metal3 ;
  RECT 645.820 165.760 649.360 166.880 ;
  LAYER metal2 ;
  RECT 645.820 165.760 649.360 166.880 ;
  LAYER metal1 ;
  RECT 645.820 165.760 649.360 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 637.140 165.760 640.680 166.880 ;
  LAYER metal3 ;
  RECT 637.140 165.760 640.680 166.880 ;
  LAYER metal2 ;
  RECT 637.140 165.760 640.680 166.880 ;
  LAYER metal1 ;
  RECT 637.140 165.760 640.680 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 628.460 165.760 632.000 166.880 ;
  LAYER metal3 ;
  RECT 628.460 165.760 632.000 166.880 ;
  LAYER metal2 ;
  RECT 628.460 165.760 632.000 166.880 ;
  LAYER metal1 ;
  RECT 628.460 165.760 632.000 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 619.780 165.760 623.320 166.880 ;
  LAYER metal3 ;
  RECT 619.780 165.760 623.320 166.880 ;
  LAYER metal2 ;
  RECT 619.780 165.760 623.320 166.880 ;
  LAYER metal1 ;
  RECT 619.780 165.760 623.320 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 576.380 165.760 579.920 166.880 ;
  LAYER metal3 ;
  RECT 576.380 165.760 579.920 166.880 ;
  LAYER metal2 ;
  RECT 576.380 165.760 579.920 166.880 ;
  LAYER metal1 ;
  RECT 576.380 165.760 579.920 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 567.700 165.760 571.240 166.880 ;
  LAYER metal3 ;
  RECT 567.700 165.760 571.240 166.880 ;
  LAYER metal2 ;
  RECT 567.700 165.760 571.240 166.880 ;
  LAYER metal1 ;
  RECT 567.700 165.760 571.240 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 559.020 165.760 562.560 166.880 ;
  LAYER metal3 ;
  RECT 559.020 165.760 562.560 166.880 ;
  LAYER metal2 ;
  RECT 559.020 165.760 562.560 166.880 ;
  LAYER metal1 ;
  RECT 559.020 165.760 562.560 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 550.340 165.760 553.880 166.880 ;
  LAYER metal3 ;
  RECT 550.340 165.760 553.880 166.880 ;
  LAYER metal2 ;
  RECT 550.340 165.760 553.880 166.880 ;
  LAYER metal1 ;
  RECT 550.340 165.760 553.880 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 541.660 165.760 545.200 166.880 ;
  LAYER metal3 ;
  RECT 541.660 165.760 545.200 166.880 ;
  LAYER metal2 ;
  RECT 541.660 165.760 545.200 166.880 ;
  LAYER metal1 ;
  RECT 541.660 165.760 545.200 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 532.980 165.760 536.520 166.880 ;
  LAYER metal3 ;
  RECT 532.980 165.760 536.520 166.880 ;
  LAYER metal2 ;
  RECT 532.980 165.760 536.520 166.880 ;
  LAYER metal1 ;
  RECT 532.980 165.760 536.520 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 489.580 165.760 493.120 166.880 ;
  LAYER metal3 ;
  RECT 489.580 165.760 493.120 166.880 ;
  LAYER metal2 ;
  RECT 489.580 165.760 493.120 166.880 ;
  LAYER metal1 ;
  RECT 489.580 165.760 493.120 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 480.900 165.760 484.440 166.880 ;
  LAYER metal3 ;
  RECT 480.900 165.760 484.440 166.880 ;
  LAYER metal2 ;
  RECT 480.900 165.760 484.440 166.880 ;
  LAYER metal1 ;
  RECT 480.900 165.760 484.440 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 472.220 165.760 475.760 166.880 ;
  LAYER metal3 ;
  RECT 472.220 165.760 475.760 166.880 ;
  LAYER metal2 ;
  RECT 472.220 165.760 475.760 166.880 ;
  LAYER metal1 ;
  RECT 472.220 165.760 475.760 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 463.540 165.760 467.080 166.880 ;
  LAYER metal3 ;
  RECT 463.540 165.760 467.080 166.880 ;
  LAYER metal2 ;
  RECT 463.540 165.760 467.080 166.880 ;
  LAYER metal1 ;
  RECT 463.540 165.760 467.080 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 454.860 165.760 458.400 166.880 ;
  LAYER metal3 ;
  RECT 454.860 165.760 458.400 166.880 ;
  LAYER metal2 ;
  RECT 454.860 165.760 458.400 166.880 ;
  LAYER metal1 ;
  RECT 454.860 165.760 458.400 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 446.180 165.760 449.720 166.880 ;
  LAYER metal3 ;
  RECT 446.180 165.760 449.720 166.880 ;
  LAYER metal2 ;
  RECT 446.180 165.760 449.720 166.880 ;
  LAYER metal1 ;
  RECT 446.180 165.760 449.720 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 402.780 165.760 406.320 166.880 ;
  LAYER metal3 ;
  RECT 402.780 165.760 406.320 166.880 ;
  LAYER metal2 ;
  RECT 402.780 165.760 406.320 166.880 ;
  LAYER metal1 ;
  RECT 402.780 165.760 406.320 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 394.100 165.760 397.640 166.880 ;
  LAYER metal3 ;
  RECT 394.100 165.760 397.640 166.880 ;
  LAYER metal2 ;
  RECT 394.100 165.760 397.640 166.880 ;
  LAYER metal1 ;
  RECT 394.100 165.760 397.640 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 385.420 165.760 388.960 166.880 ;
  LAYER metal3 ;
  RECT 385.420 165.760 388.960 166.880 ;
  LAYER metal2 ;
  RECT 385.420 165.760 388.960 166.880 ;
  LAYER metal1 ;
  RECT 385.420 165.760 388.960 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 376.740 165.760 380.280 166.880 ;
  LAYER metal3 ;
  RECT 376.740 165.760 380.280 166.880 ;
  LAYER metal2 ;
  RECT 376.740 165.760 380.280 166.880 ;
  LAYER metal1 ;
  RECT 376.740 165.760 380.280 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 368.060 165.760 371.600 166.880 ;
  LAYER metal3 ;
  RECT 368.060 165.760 371.600 166.880 ;
  LAYER metal2 ;
  RECT 368.060 165.760 371.600 166.880 ;
  LAYER metal1 ;
  RECT 368.060 165.760 371.600 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 359.380 165.760 362.920 166.880 ;
  LAYER metal3 ;
  RECT 359.380 165.760 362.920 166.880 ;
  LAYER metal2 ;
  RECT 359.380 165.760 362.920 166.880 ;
  LAYER metal1 ;
  RECT 359.380 165.760 362.920 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.980 165.760 319.520 166.880 ;
  LAYER metal3 ;
  RECT 315.980 165.760 319.520 166.880 ;
  LAYER metal2 ;
  RECT 315.980 165.760 319.520 166.880 ;
  LAYER metal1 ;
  RECT 315.980 165.760 319.520 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 307.300 165.760 310.840 166.880 ;
  LAYER metal3 ;
  RECT 307.300 165.760 310.840 166.880 ;
  LAYER metal2 ;
  RECT 307.300 165.760 310.840 166.880 ;
  LAYER metal1 ;
  RECT 307.300 165.760 310.840 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 298.620 165.760 302.160 166.880 ;
  LAYER metal3 ;
  RECT 298.620 165.760 302.160 166.880 ;
  LAYER metal2 ;
  RECT 298.620 165.760 302.160 166.880 ;
  LAYER metal1 ;
  RECT 298.620 165.760 302.160 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 289.940 165.760 293.480 166.880 ;
  LAYER metal3 ;
  RECT 289.940 165.760 293.480 166.880 ;
  LAYER metal2 ;
  RECT 289.940 165.760 293.480 166.880 ;
  LAYER metal1 ;
  RECT 289.940 165.760 293.480 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 281.260 165.760 284.800 166.880 ;
  LAYER metal3 ;
  RECT 281.260 165.760 284.800 166.880 ;
  LAYER metal2 ;
  RECT 281.260 165.760 284.800 166.880 ;
  LAYER metal1 ;
  RECT 281.260 165.760 284.800 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 272.580 165.760 276.120 166.880 ;
  LAYER metal3 ;
  RECT 272.580 165.760 276.120 166.880 ;
  LAYER metal2 ;
  RECT 272.580 165.760 276.120 166.880 ;
  LAYER metal1 ;
  RECT 272.580 165.760 276.120 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 229.180 165.760 232.720 166.880 ;
  LAYER metal3 ;
  RECT 229.180 165.760 232.720 166.880 ;
  LAYER metal2 ;
  RECT 229.180 165.760 232.720 166.880 ;
  LAYER metal1 ;
  RECT 229.180 165.760 232.720 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 220.500 165.760 224.040 166.880 ;
  LAYER metal3 ;
  RECT 220.500 165.760 224.040 166.880 ;
  LAYER metal2 ;
  RECT 220.500 165.760 224.040 166.880 ;
  LAYER metal1 ;
  RECT 220.500 165.760 224.040 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 211.820 165.760 215.360 166.880 ;
  LAYER metal3 ;
  RECT 211.820 165.760 215.360 166.880 ;
  LAYER metal2 ;
  RECT 211.820 165.760 215.360 166.880 ;
  LAYER metal1 ;
  RECT 211.820 165.760 215.360 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 203.140 165.760 206.680 166.880 ;
  LAYER metal3 ;
  RECT 203.140 165.760 206.680 166.880 ;
  LAYER metal2 ;
  RECT 203.140 165.760 206.680 166.880 ;
  LAYER metal1 ;
  RECT 203.140 165.760 206.680 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 194.460 165.760 198.000 166.880 ;
  LAYER metal3 ;
  RECT 194.460 165.760 198.000 166.880 ;
  LAYER metal2 ;
  RECT 194.460 165.760 198.000 166.880 ;
  LAYER metal1 ;
  RECT 194.460 165.760 198.000 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 185.780 165.760 189.320 166.880 ;
  LAYER metal3 ;
  RECT 185.780 165.760 189.320 166.880 ;
  LAYER metal2 ;
  RECT 185.780 165.760 189.320 166.880 ;
  LAYER metal1 ;
  RECT 185.780 165.760 189.320 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 142.380 165.760 145.920 166.880 ;
  LAYER metal3 ;
  RECT 142.380 165.760 145.920 166.880 ;
  LAYER metal2 ;
  RECT 142.380 165.760 145.920 166.880 ;
  LAYER metal1 ;
  RECT 142.380 165.760 145.920 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 133.700 165.760 137.240 166.880 ;
  LAYER metal3 ;
  RECT 133.700 165.760 137.240 166.880 ;
  LAYER metal2 ;
  RECT 133.700 165.760 137.240 166.880 ;
  LAYER metal1 ;
  RECT 133.700 165.760 137.240 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 125.020 165.760 128.560 166.880 ;
  LAYER metal3 ;
  RECT 125.020 165.760 128.560 166.880 ;
  LAYER metal2 ;
  RECT 125.020 165.760 128.560 166.880 ;
  LAYER metal1 ;
  RECT 125.020 165.760 128.560 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 116.340 165.760 119.880 166.880 ;
  LAYER metal3 ;
  RECT 116.340 165.760 119.880 166.880 ;
  LAYER metal2 ;
  RECT 116.340 165.760 119.880 166.880 ;
  LAYER metal1 ;
  RECT 116.340 165.760 119.880 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 107.660 165.760 111.200 166.880 ;
  LAYER metal3 ;
  RECT 107.660 165.760 111.200 166.880 ;
  LAYER metal2 ;
  RECT 107.660 165.760 111.200 166.880 ;
  LAYER metal1 ;
  RECT 107.660 165.760 111.200 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 98.980 165.760 102.520 166.880 ;
  LAYER metal3 ;
  RECT 98.980 165.760 102.520 166.880 ;
  LAYER metal2 ;
  RECT 98.980 165.760 102.520 166.880 ;
  LAYER metal1 ;
  RECT 98.980 165.760 102.520 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 55.580 165.760 59.120 166.880 ;
  LAYER metal3 ;
  RECT 55.580 165.760 59.120 166.880 ;
  LAYER metal2 ;
  RECT 55.580 165.760 59.120 166.880 ;
  LAYER metal1 ;
  RECT 55.580 165.760 59.120 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 46.900 165.760 50.440 166.880 ;
  LAYER metal3 ;
  RECT 46.900 165.760 50.440 166.880 ;
  LAYER metal2 ;
  RECT 46.900 165.760 50.440 166.880 ;
  LAYER metal1 ;
  RECT 46.900 165.760 50.440 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 38.220 165.760 41.760 166.880 ;
  LAYER metal3 ;
  RECT 38.220 165.760 41.760 166.880 ;
  LAYER metal2 ;
  RECT 38.220 165.760 41.760 166.880 ;
  LAYER metal1 ;
  RECT 38.220 165.760 41.760 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 29.540 165.760 33.080 166.880 ;
  LAYER metal3 ;
  RECT 29.540 165.760 33.080 166.880 ;
  LAYER metal2 ;
  RECT 29.540 165.760 33.080 166.880 ;
  LAYER metal1 ;
  RECT 29.540 165.760 33.080 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 20.860 165.760 24.400 166.880 ;
  LAYER metal3 ;
  RECT 20.860 165.760 24.400 166.880 ;
  LAYER metal2 ;
  RECT 20.860 165.760 24.400 166.880 ;
  LAYER metal1 ;
  RECT 20.860 165.760 24.400 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 12.180 165.760 15.720 166.880 ;
  LAYER metal3 ;
  RECT 12.180 165.760 15.720 166.880 ;
  LAYER metal2 ;
  RECT 12.180 165.760 15.720 166.880 ;
  LAYER metal1 ;
  RECT 12.180 165.760 15.720 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1857.300 0.000 1860.840 1.120 ;
  LAYER metal3 ;
  RECT 1857.300 0.000 1860.840 1.120 ;
  LAYER metal2 ;
  RECT 1857.300 0.000 1860.840 1.120 ;
  LAYER metal1 ;
  RECT 1857.300 0.000 1860.840 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1848.620 0.000 1852.160 1.120 ;
  LAYER metal3 ;
  RECT 1848.620 0.000 1852.160 1.120 ;
  LAYER metal2 ;
  RECT 1848.620 0.000 1852.160 1.120 ;
  LAYER metal1 ;
  RECT 1848.620 0.000 1852.160 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1839.940 0.000 1843.480 1.120 ;
  LAYER metal3 ;
  RECT 1839.940 0.000 1843.480 1.120 ;
  LAYER metal2 ;
  RECT 1839.940 0.000 1843.480 1.120 ;
  LAYER metal1 ;
  RECT 1839.940 0.000 1843.480 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1831.260 0.000 1834.800 1.120 ;
  LAYER metal3 ;
  RECT 1831.260 0.000 1834.800 1.120 ;
  LAYER metal2 ;
  RECT 1831.260 0.000 1834.800 1.120 ;
  LAYER metal1 ;
  RECT 1831.260 0.000 1834.800 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1822.580 0.000 1826.120 1.120 ;
  LAYER metal3 ;
  RECT 1822.580 0.000 1826.120 1.120 ;
  LAYER metal2 ;
  RECT 1822.580 0.000 1826.120 1.120 ;
  LAYER metal1 ;
  RECT 1822.580 0.000 1826.120 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1813.900 0.000 1817.440 1.120 ;
  LAYER metal3 ;
  RECT 1813.900 0.000 1817.440 1.120 ;
  LAYER metal2 ;
  RECT 1813.900 0.000 1817.440 1.120 ;
  LAYER metal1 ;
  RECT 1813.900 0.000 1817.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1753.140 0.000 1756.680 1.120 ;
  LAYER metal3 ;
  RECT 1753.140 0.000 1756.680 1.120 ;
  LAYER metal2 ;
  RECT 1753.140 0.000 1756.680 1.120 ;
  LAYER metal1 ;
  RECT 1753.140 0.000 1756.680 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1744.460 0.000 1748.000 1.120 ;
  LAYER metal3 ;
  RECT 1744.460 0.000 1748.000 1.120 ;
  LAYER metal2 ;
  RECT 1744.460 0.000 1748.000 1.120 ;
  LAYER metal1 ;
  RECT 1744.460 0.000 1748.000 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1735.780 0.000 1739.320 1.120 ;
  LAYER metal3 ;
  RECT 1735.780 0.000 1739.320 1.120 ;
  LAYER metal2 ;
  RECT 1735.780 0.000 1739.320 1.120 ;
  LAYER metal1 ;
  RECT 1735.780 0.000 1739.320 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1727.100 0.000 1730.640 1.120 ;
  LAYER metal3 ;
  RECT 1727.100 0.000 1730.640 1.120 ;
  LAYER metal2 ;
  RECT 1727.100 0.000 1730.640 1.120 ;
  LAYER metal1 ;
  RECT 1727.100 0.000 1730.640 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1718.420 0.000 1721.960 1.120 ;
  LAYER metal3 ;
  RECT 1718.420 0.000 1721.960 1.120 ;
  LAYER metal2 ;
  RECT 1718.420 0.000 1721.960 1.120 ;
  LAYER metal1 ;
  RECT 1718.420 0.000 1721.960 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1709.740 0.000 1713.280 1.120 ;
  LAYER metal3 ;
  RECT 1709.740 0.000 1713.280 1.120 ;
  LAYER metal2 ;
  RECT 1709.740 0.000 1713.280 1.120 ;
  LAYER metal1 ;
  RECT 1709.740 0.000 1713.280 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1648.980 0.000 1652.520 1.120 ;
  LAYER metal3 ;
  RECT 1648.980 0.000 1652.520 1.120 ;
  LAYER metal2 ;
  RECT 1648.980 0.000 1652.520 1.120 ;
  LAYER metal1 ;
  RECT 1648.980 0.000 1652.520 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1640.300 0.000 1643.840 1.120 ;
  LAYER metal3 ;
  RECT 1640.300 0.000 1643.840 1.120 ;
  LAYER metal2 ;
  RECT 1640.300 0.000 1643.840 1.120 ;
  LAYER metal1 ;
  RECT 1640.300 0.000 1643.840 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1631.620 0.000 1635.160 1.120 ;
  LAYER metal3 ;
  RECT 1631.620 0.000 1635.160 1.120 ;
  LAYER metal2 ;
  RECT 1631.620 0.000 1635.160 1.120 ;
  LAYER metal1 ;
  RECT 1631.620 0.000 1635.160 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1622.940 0.000 1626.480 1.120 ;
  LAYER metal3 ;
  RECT 1622.940 0.000 1626.480 1.120 ;
  LAYER metal2 ;
  RECT 1622.940 0.000 1626.480 1.120 ;
  LAYER metal1 ;
  RECT 1622.940 0.000 1626.480 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1614.260 0.000 1617.800 1.120 ;
  LAYER metal3 ;
  RECT 1614.260 0.000 1617.800 1.120 ;
  LAYER metal2 ;
  RECT 1614.260 0.000 1617.800 1.120 ;
  LAYER metal1 ;
  RECT 1614.260 0.000 1617.800 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1605.580 0.000 1609.120 1.120 ;
  LAYER metal3 ;
  RECT 1605.580 0.000 1609.120 1.120 ;
  LAYER metal2 ;
  RECT 1605.580 0.000 1609.120 1.120 ;
  LAYER metal1 ;
  RECT 1605.580 0.000 1609.120 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1544.200 0.000 1547.740 1.120 ;
  LAYER metal3 ;
  RECT 1544.200 0.000 1547.740 1.120 ;
  LAYER metal2 ;
  RECT 1544.200 0.000 1547.740 1.120 ;
  LAYER metal1 ;
  RECT 1544.200 0.000 1547.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1535.520 0.000 1539.060 1.120 ;
  LAYER metal3 ;
  RECT 1535.520 0.000 1539.060 1.120 ;
  LAYER metal2 ;
  RECT 1535.520 0.000 1539.060 1.120 ;
  LAYER metal1 ;
  RECT 1535.520 0.000 1539.060 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1526.840 0.000 1530.380 1.120 ;
  LAYER metal3 ;
  RECT 1526.840 0.000 1530.380 1.120 ;
  LAYER metal2 ;
  RECT 1526.840 0.000 1530.380 1.120 ;
  LAYER metal1 ;
  RECT 1526.840 0.000 1530.380 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1518.160 0.000 1521.700 1.120 ;
  LAYER metal3 ;
  RECT 1518.160 0.000 1521.700 1.120 ;
  LAYER metal2 ;
  RECT 1518.160 0.000 1521.700 1.120 ;
  LAYER metal1 ;
  RECT 1518.160 0.000 1521.700 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1509.480 0.000 1513.020 1.120 ;
  LAYER metal3 ;
  RECT 1509.480 0.000 1513.020 1.120 ;
  LAYER metal2 ;
  RECT 1509.480 0.000 1513.020 1.120 ;
  LAYER metal1 ;
  RECT 1509.480 0.000 1513.020 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1500.800 0.000 1504.340 1.120 ;
  LAYER metal3 ;
  RECT 1500.800 0.000 1504.340 1.120 ;
  LAYER metal2 ;
  RECT 1500.800 0.000 1504.340 1.120 ;
  LAYER metal1 ;
  RECT 1500.800 0.000 1504.340 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1453.680 0.000 1457.220 1.120 ;
  LAYER metal3 ;
  RECT 1453.680 0.000 1457.220 1.120 ;
  LAYER metal2 ;
  RECT 1453.680 0.000 1457.220 1.120 ;
  LAYER metal1 ;
  RECT 1453.680 0.000 1457.220 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1431.360 0.000 1434.900 1.120 ;
  LAYER metal3 ;
  RECT 1431.360 0.000 1434.900 1.120 ;
  LAYER metal2 ;
  RECT 1431.360 0.000 1434.900 1.120 ;
  LAYER metal1 ;
  RECT 1431.360 0.000 1434.900 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1422.680 0.000 1426.220 1.120 ;
  LAYER metal3 ;
  RECT 1422.680 0.000 1426.220 1.120 ;
  LAYER metal2 ;
  RECT 1422.680 0.000 1426.220 1.120 ;
  LAYER metal1 ;
  RECT 1422.680 0.000 1426.220 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1414.000 0.000 1417.540 1.120 ;
  LAYER metal3 ;
  RECT 1414.000 0.000 1417.540 1.120 ;
  LAYER metal2 ;
  RECT 1414.000 0.000 1417.540 1.120 ;
  LAYER metal1 ;
  RECT 1414.000 0.000 1417.540 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1405.320 0.000 1408.860 1.120 ;
  LAYER metal3 ;
  RECT 1405.320 0.000 1408.860 1.120 ;
  LAYER metal2 ;
  RECT 1405.320 0.000 1408.860 1.120 ;
  LAYER metal1 ;
  RECT 1405.320 0.000 1408.860 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1396.640 0.000 1400.180 1.120 ;
  LAYER metal3 ;
  RECT 1396.640 0.000 1400.180 1.120 ;
  LAYER metal2 ;
  RECT 1396.640 0.000 1400.180 1.120 ;
  LAYER metal1 ;
  RECT 1396.640 0.000 1400.180 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1353.240 0.000 1356.780 1.120 ;
  LAYER metal3 ;
  RECT 1353.240 0.000 1356.780 1.120 ;
  LAYER metal2 ;
  RECT 1353.240 0.000 1356.780 1.120 ;
  LAYER metal1 ;
  RECT 1353.240 0.000 1356.780 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1340.220 0.000 1343.760 1.120 ;
  LAYER metal3 ;
  RECT 1340.220 0.000 1343.760 1.120 ;
  LAYER metal2 ;
  RECT 1340.220 0.000 1343.760 1.120 ;
  LAYER metal1 ;
  RECT 1340.220 0.000 1343.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1318.520 0.000 1322.060 1.120 ;
  LAYER metal3 ;
  RECT 1318.520 0.000 1322.060 1.120 ;
  LAYER metal2 ;
  RECT 1318.520 0.000 1322.060 1.120 ;
  LAYER metal1 ;
  RECT 1318.520 0.000 1322.060 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1309.840 0.000 1313.380 1.120 ;
  LAYER metal3 ;
  RECT 1309.840 0.000 1313.380 1.120 ;
  LAYER metal2 ;
  RECT 1309.840 0.000 1313.380 1.120 ;
  LAYER metal1 ;
  RECT 1309.840 0.000 1313.380 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1301.160 0.000 1304.700 1.120 ;
  LAYER metal3 ;
  RECT 1301.160 0.000 1304.700 1.120 ;
  LAYER metal2 ;
  RECT 1301.160 0.000 1304.700 1.120 ;
  LAYER metal1 ;
  RECT 1301.160 0.000 1304.700 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1292.480 0.000 1296.020 1.120 ;
  LAYER metal3 ;
  RECT 1292.480 0.000 1296.020 1.120 ;
  LAYER metal2 ;
  RECT 1292.480 0.000 1296.020 1.120 ;
  LAYER metal1 ;
  RECT 1292.480 0.000 1296.020 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1249.080 0.000 1252.620 1.120 ;
  LAYER metal3 ;
  RECT 1249.080 0.000 1252.620 1.120 ;
  LAYER metal2 ;
  RECT 1249.080 0.000 1252.620 1.120 ;
  LAYER metal1 ;
  RECT 1249.080 0.000 1252.620 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1240.400 0.000 1243.940 1.120 ;
  LAYER metal3 ;
  RECT 1240.400 0.000 1243.940 1.120 ;
  LAYER metal2 ;
  RECT 1240.400 0.000 1243.940 1.120 ;
  LAYER metal1 ;
  RECT 1240.400 0.000 1243.940 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1227.380 0.000 1230.920 1.120 ;
  LAYER metal3 ;
  RECT 1227.380 0.000 1230.920 1.120 ;
  LAYER metal2 ;
  RECT 1227.380 0.000 1230.920 1.120 ;
  LAYER metal1 ;
  RECT 1227.380 0.000 1230.920 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1205.060 0.000 1208.600 1.120 ;
  LAYER metal3 ;
  RECT 1205.060 0.000 1208.600 1.120 ;
  LAYER metal2 ;
  RECT 1205.060 0.000 1208.600 1.120 ;
  LAYER metal1 ;
  RECT 1205.060 0.000 1208.600 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1196.380 0.000 1199.920 1.120 ;
  LAYER metal3 ;
  RECT 1196.380 0.000 1199.920 1.120 ;
  LAYER metal2 ;
  RECT 1196.380 0.000 1199.920 1.120 ;
  LAYER metal1 ;
  RECT 1196.380 0.000 1199.920 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1187.700 0.000 1191.240 1.120 ;
  LAYER metal3 ;
  RECT 1187.700 0.000 1191.240 1.120 ;
  LAYER metal2 ;
  RECT 1187.700 0.000 1191.240 1.120 ;
  LAYER metal1 ;
  RECT 1187.700 0.000 1191.240 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1144.300 0.000 1147.840 1.120 ;
  LAYER metal3 ;
  RECT 1144.300 0.000 1147.840 1.120 ;
  LAYER metal2 ;
  RECT 1144.300 0.000 1147.840 1.120 ;
  LAYER metal1 ;
  RECT 1144.300 0.000 1147.840 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1135.620 0.000 1139.160 1.120 ;
  LAYER metal3 ;
  RECT 1135.620 0.000 1139.160 1.120 ;
  LAYER metal2 ;
  RECT 1135.620 0.000 1139.160 1.120 ;
  LAYER metal1 ;
  RECT 1135.620 0.000 1139.160 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1126.940 0.000 1130.480 1.120 ;
  LAYER metal3 ;
  RECT 1126.940 0.000 1130.480 1.120 ;
  LAYER metal2 ;
  RECT 1126.940 0.000 1130.480 1.120 ;
  LAYER metal1 ;
  RECT 1126.940 0.000 1130.480 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1114.540 0.000 1118.080 1.120 ;
  LAYER metal3 ;
  RECT 1114.540 0.000 1118.080 1.120 ;
  LAYER metal2 ;
  RECT 1114.540 0.000 1118.080 1.120 ;
  LAYER metal1 ;
  RECT 1114.540 0.000 1118.080 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1092.220 0.000 1095.760 1.120 ;
  LAYER metal3 ;
  RECT 1092.220 0.000 1095.760 1.120 ;
  LAYER metal2 ;
  RECT 1092.220 0.000 1095.760 1.120 ;
  LAYER metal1 ;
  RECT 1092.220 0.000 1095.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1083.540 0.000 1087.080 1.120 ;
  LAYER metal3 ;
  RECT 1083.540 0.000 1087.080 1.120 ;
  LAYER metal2 ;
  RECT 1083.540 0.000 1087.080 1.120 ;
  LAYER metal1 ;
  RECT 1083.540 0.000 1087.080 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1040.140 0.000 1043.680 1.120 ;
  LAYER metal3 ;
  RECT 1040.140 0.000 1043.680 1.120 ;
  LAYER metal2 ;
  RECT 1040.140 0.000 1043.680 1.120 ;
  LAYER metal1 ;
  RECT 1040.140 0.000 1043.680 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1031.460 0.000 1035.000 1.120 ;
  LAYER metal3 ;
  RECT 1031.460 0.000 1035.000 1.120 ;
  LAYER metal2 ;
  RECT 1031.460 0.000 1035.000 1.120 ;
  LAYER metal1 ;
  RECT 1031.460 0.000 1035.000 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1022.780 0.000 1026.320 1.120 ;
  LAYER metal3 ;
  RECT 1022.780 0.000 1026.320 1.120 ;
  LAYER metal2 ;
  RECT 1022.780 0.000 1026.320 1.120 ;
  LAYER metal1 ;
  RECT 1022.780 0.000 1026.320 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1014.100 0.000 1017.640 1.120 ;
  LAYER metal3 ;
  RECT 1014.100 0.000 1017.640 1.120 ;
  LAYER metal2 ;
  RECT 1014.100 0.000 1017.640 1.120 ;
  LAYER metal1 ;
  RECT 1014.100 0.000 1017.640 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1001.080 0.000 1004.620 1.120 ;
  LAYER metal3 ;
  RECT 1001.080 0.000 1004.620 1.120 ;
  LAYER metal2 ;
  RECT 1001.080 0.000 1004.620 1.120 ;
  LAYER metal1 ;
  RECT 1001.080 0.000 1004.620 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 965.120 0.000 968.660 1.120 ;
  LAYER metal3 ;
  RECT 965.120 0.000 968.660 1.120 ;
  LAYER metal2 ;
  RECT 965.120 0.000 968.660 1.120 ;
  LAYER metal1 ;
  RECT 965.120 0.000 968.660 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 891.960 0.000 895.500 1.120 ;
  LAYER metal3 ;
  RECT 891.960 0.000 895.500 1.120 ;
  LAYER metal2 ;
  RECT 891.960 0.000 895.500 1.120 ;
  LAYER metal1 ;
  RECT 891.960 0.000 895.500 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 883.280 0.000 886.820 1.120 ;
  LAYER metal3 ;
  RECT 883.280 0.000 886.820 1.120 ;
  LAYER metal2 ;
  RECT 883.280 0.000 886.820 1.120 ;
  LAYER metal1 ;
  RECT 883.280 0.000 886.820 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 874.600 0.000 878.140 1.120 ;
  LAYER metal3 ;
  RECT 874.600 0.000 878.140 1.120 ;
  LAYER metal2 ;
  RECT 874.600 0.000 878.140 1.120 ;
  LAYER metal1 ;
  RECT 874.600 0.000 878.140 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 865.920 0.000 869.460 1.120 ;
  LAYER metal3 ;
  RECT 865.920 0.000 869.460 1.120 ;
  LAYER metal2 ;
  RECT 865.920 0.000 869.460 1.120 ;
  LAYER metal1 ;
  RECT 865.920 0.000 869.460 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 857.240 0.000 860.780 1.120 ;
  LAYER metal3 ;
  RECT 857.240 0.000 860.780 1.120 ;
  LAYER metal2 ;
  RECT 857.240 0.000 860.780 1.120 ;
  LAYER metal1 ;
  RECT 857.240 0.000 860.780 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 848.560 0.000 852.100 1.120 ;
  LAYER metal3 ;
  RECT 848.560 0.000 852.100 1.120 ;
  LAYER metal2 ;
  RECT 848.560 0.000 852.100 1.120 ;
  LAYER metal1 ;
  RECT 848.560 0.000 852.100 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 787.800 0.000 791.340 1.120 ;
  LAYER metal3 ;
  RECT 787.800 0.000 791.340 1.120 ;
  LAYER metal2 ;
  RECT 787.800 0.000 791.340 1.120 ;
  LAYER metal1 ;
  RECT 787.800 0.000 791.340 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 779.120 0.000 782.660 1.120 ;
  LAYER metal3 ;
  RECT 779.120 0.000 782.660 1.120 ;
  LAYER metal2 ;
  RECT 779.120 0.000 782.660 1.120 ;
  LAYER metal1 ;
  RECT 779.120 0.000 782.660 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 770.440 0.000 773.980 1.120 ;
  LAYER metal3 ;
  RECT 770.440 0.000 773.980 1.120 ;
  LAYER metal2 ;
  RECT 770.440 0.000 773.980 1.120 ;
  LAYER metal1 ;
  RECT 770.440 0.000 773.980 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 761.760 0.000 765.300 1.120 ;
  LAYER metal3 ;
  RECT 761.760 0.000 765.300 1.120 ;
  LAYER metal2 ;
  RECT 761.760 0.000 765.300 1.120 ;
  LAYER metal1 ;
  RECT 761.760 0.000 765.300 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 753.080 0.000 756.620 1.120 ;
  LAYER metal3 ;
  RECT 753.080 0.000 756.620 1.120 ;
  LAYER metal2 ;
  RECT 753.080 0.000 756.620 1.120 ;
  LAYER metal1 ;
  RECT 753.080 0.000 756.620 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 744.400 0.000 747.940 1.120 ;
  LAYER metal3 ;
  RECT 744.400 0.000 747.940 1.120 ;
  LAYER metal2 ;
  RECT 744.400 0.000 747.940 1.120 ;
  LAYER metal1 ;
  RECT 744.400 0.000 747.940 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 683.020 0.000 686.560 1.120 ;
  LAYER metal3 ;
  RECT 683.020 0.000 686.560 1.120 ;
  LAYER metal2 ;
  RECT 683.020 0.000 686.560 1.120 ;
  LAYER metal1 ;
  RECT 683.020 0.000 686.560 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 674.340 0.000 677.880 1.120 ;
  LAYER metal3 ;
  RECT 674.340 0.000 677.880 1.120 ;
  LAYER metal2 ;
  RECT 674.340 0.000 677.880 1.120 ;
  LAYER metal1 ;
  RECT 674.340 0.000 677.880 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 665.660 0.000 669.200 1.120 ;
  LAYER metal3 ;
  RECT 665.660 0.000 669.200 1.120 ;
  LAYER metal2 ;
  RECT 665.660 0.000 669.200 1.120 ;
  LAYER metal1 ;
  RECT 665.660 0.000 669.200 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 656.980 0.000 660.520 1.120 ;
  LAYER metal3 ;
  RECT 656.980 0.000 660.520 1.120 ;
  LAYER metal2 ;
  RECT 656.980 0.000 660.520 1.120 ;
  LAYER metal1 ;
  RECT 656.980 0.000 660.520 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 648.300 0.000 651.840 1.120 ;
  LAYER metal3 ;
  RECT 648.300 0.000 651.840 1.120 ;
  LAYER metal2 ;
  RECT 648.300 0.000 651.840 1.120 ;
  LAYER metal1 ;
  RECT 648.300 0.000 651.840 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 639.620 0.000 643.160 1.120 ;
  LAYER metal3 ;
  RECT 639.620 0.000 643.160 1.120 ;
  LAYER metal2 ;
  RECT 639.620 0.000 643.160 1.120 ;
  LAYER metal1 ;
  RECT 639.620 0.000 643.160 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 592.500 0.000 596.040 1.120 ;
  LAYER metal3 ;
  RECT 592.500 0.000 596.040 1.120 ;
  LAYER metal2 ;
  RECT 592.500 0.000 596.040 1.120 ;
  LAYER metal1 ;
  RECT 592.500 0.000 596.040 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal3 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal2 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal1 ;
  RECT 570.180 0.000 573.720 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 561.500 0.000 565.040 1.120 ;
  LAYER metal3 ;
  RECT 561.500 0.000 565.040 1.120 ;
  LAYER metal2 ;
  RECT 561.500 0.000 565.040 1.120 ;
  LAYER metal1 ;
  RECT 561.500 0.000 565.040 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 552.820 0.000 556.360 1.120 ;
  LAYER metal3 ;
  RECT 552.820 0.000 556.360 1.120 ;
  LAYER metal2 ;
  RECT 552.820 0.000 556.360 1.120 ;
  LAYER metal1 ;
  RECT 552.820 0.000 556.360 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 544.140 0.000 547.680 1.120 ;
  LAYER metal3 ;
  RECT 544.140 0.000 547.680 1.120 ;
  LAYER metal2 ;
  RECT 544.140 0.000 547.680 1.120 ;
  LAYER metal1 ;
  RECT 544.140 0.000 547.680 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 535.460 0.000 539.000 1.120 ;
  LAYER metal3 ;
  RECT 535.460 0.000 539.000 1.120 ;
  LAYER metal2 ;
  RECT 535.460 0.000 539.000 1.120 ;
  LAYER metal1 ;
  RECT 535.460 0.000 539.000 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 492.060 0.000 495.600 1.120 ;
  LAYER metal3 ;
  RECT 492.060 0.000 495.600 1.120 ;
  LAYER metal2 ;
  RECT 492.060 0.000 495.600 1.120 ;
  LAYER metal1 ;
  RECT 492.060 0.000 495.600 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 479.040 0.000 482.580 1.120 ;
  LAYER metal3 ;
  RECT 479.040 0.000 482.580 1.120 ;
  LAYER metal2 ;
  RECT 479.040 0.000 482.580 1.120 ;
  LAYER metal1 ;
  RECT 479.040 0.000 482.580 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 457.340 0.000 460.880 1.120 ;
  LAYER metal3 ;
  RECT 457.340 0.000 460.880 1.120 ;
  LAYER metal2 ;
  RECT 457.340 0.000 460.880 1.120 ;
  LAYER metal1 ;
  RECT 457.340 0.000 460.880 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 448.660 0.000 452.200 1.120 ;
  LAYER metal3 ;
  RECT 448.660 0.000 452.200 1.120 ;
  LAYER metal2 ;
  RECT 448.660 0.000 452.200 1.120 ;
  LAYER metal1 ;
  RECT 448.660 0.000 452.200 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 439.980 0.000 443.520 1.120 ;
  LAYER metal3 ;
  RECT 439.980 0.000 443.520 1.120 ;
  LAYER metal2 ;
  RECT 439.980 0.000 443.520 1.120 ;
  LAYER metal1 ;
  RECT 439.980 0.000 443.520 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER metal3 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER metal2 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER metal1 ;
  RECT 431.300 0.000 434.840 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 387.900 0.000 391.440 1.120 ;
  LAYER metal3 ;
  RECT 387.900 0.000 391.440 1.120 ;
  LAYER metal2 ;
  RECT 387.900 0.000 391.440 1.120 ;
  LAYER metal1 ;
  RECT 387.900 0.000 391.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 379.220 0.000 382.760 1.120 ;
  LAYER metal3 ;
  RECT 379.220 0.000 382.760 1.120 ;
  LAYER metal2 ;
  RECT 379.220 0.000 382.760 1.120 ;
  LAYER metal1 ;
  RECT 379.220 0.000 382.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 366.200 0.000 369.740 1.120 ;
  LAYER metal3 ;
  RECT 366.200 0.000 369.740 1.120 ;
  LAYER metal2 ;
  RECT 366.200 0.000 369.740 1.120 ;
  LAYER metal1 ;
  RECT 366.200 0.000 369.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 343.880 0.000 347.420 1.120 ;
  LAYER metal3 ;
  RECT 343.880 0.000 347.420 1.120 ;
  LAYER metal2 ;
  RECT 343.880 0.000 347.420 1.120 ;
  LAYER metal1 ;
  RECT 343.880 0.000 347.420 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 335.200 0.000 338.740 1.120 ;
  LAYER metal3 ;
  RECT 335.200 0.000 338.740 1.120 ;
  LAYER metal2 ;
  RECT 335.200 0.000 338.740 1.120 ;
  LAYER metal1 ;
  RECT 335.200 0.000 338.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 326.520 0.000 330.060 1.120 ;
  LAYER metal3 ;
  RECT 326.520 0.000 330.060 1.120 ;
  LAYER metal2 ;
  RECT 326.520 0.000 330.060 1.120 ;
  LAYER metal1 ;
  RECT 326.520 0.000 330.060 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER metal3 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER metal2 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER metal1 ;
  RECT 283.120 0.000 286.660 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal3 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal2 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal1 ;
  RECT 274.440 0.000 277.980 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 265.760 0.000 269.300 1.120 ;
  LAYER metal3 ;
  RECT 265.760 0.000 269.300 1.120 ;
  LAYER metal2 ;
  RECT 265.760 0.000 269.300 1.120 ;
  LAYER metal1 ;
  RECT 265.760 0.000 269.300 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER metal3 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER metal2 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER metal1 ;
  RECT 253.360 0.000 256.900 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 231.040 0.000 234.580 1.120 ;
  LAYER metal3 ;
  RECT 231.040 0.000 234.580 1.120 ;
  LAYER metal2 ;
  RECT 231.040 0.000 234.580 1.120 ;
  LAYER metal1 ;
  RECT 231.040 0.000 234.580 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 222.360 0.000 225.900 1.120 ;
  LAYER metal3 ;
  RECT 222.360 0.000 225.900 1.120 ;
  LAYER metal2 ;
  RECT 222.360 0.000 225.900 1.120 ;
  LAYER metal1 ;
  RECT 222.360 0.000 225.900 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 178.960 0.000 182.500 1.120 ;
  LAYER metal3 ;
  RECT 178.960 0.000 182.500 1.120 ;
  LAYER metal2 ;
  RECT 178.960 0.000 182.500 1.120 ;
  LAYER metal1 ;
  RECT 178.960 0.000 182.500 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 170.280 0.000 173.820 1.120 ;
  LAYER metal3 ;
  RECT 170.280 0.000 173.820 1.120 ;
  LAYER metal2 ;
  RECT 170.280 0.000 173.820 1.120 ;
  LAYER metal1 ;
  RECT 170.280 0.000 173.820 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 161.600 0.000 165.140 1.120 ;
  LAYER metal3 ;
  RECT 161.600 0.000 165.140 1.120 ;
  LAYER metal2 ;
  RECT 161.600 0.000 165.140 1.120 ;
  LAYER metal1 ;
  RECT 161.600 0.000 165.140 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 152.920 0.000 156.460 1.120 ;
  LAYER metal3 ;
  RECT 152.920 0.000 156.460 1.120 ;
  LAYER metal2 ;
  RECT 152.920 0.000 156.460 1.120 ;
  LAYER metal1 ;
  RECT 152.920 0.000 156.460 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal3 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal2 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal1 ;
  RECT 139.900 0.000 143.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 118.200 0.000 121.740 1.120 ;
  LAYER metal3 ;
  RECT 118.200 0.000 121.740 1.120 ;
  LAYER metal2 ;
  RECT 118.200 0.000 121.740 1.120 ;
  LAYER metal1 ;
  RECT 118.200 0.000 121.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 74.800 0.000 78.340 1.120 ;
  LAYER metal3 ;
  RECT 74.800 0.000 78.340 1.120 ;
  LAYER metal2 ;
  RECT 74.800 0.000 78.340 1.120 ;
  LAYER metal1 ;
  RECT 74.800 0.000 78.340 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 66.120 0.000 69.660 1.120 ;
  LAYER metal3 ;
  RECT 66.120 0.000 69.660 1.120 ;
  LAYER metal2 ;
  RECT 66.120 0.000 69.660 1.120 ;
  LAYER metal1 ;
  RECT 66.120 0.000 69.660 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 57.440 0.000 60.980 1.120 ;
  LAYER metal3 ;
  RECT 57.440 0.000 60.980 1.120 ;
  LAYER metal2 ;
  RECT 57.440 0.000 60.980 1.120 ;
  LAYER metal1 ;
  RECT 57.440 0.000 60.980 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 48.760 0.000 52.300 1.120 ;
  LAYER metal3 ;
  RECT 48.760 0.000 52.300 1.120 ;
  LAYER metal2 ;
  RECT 48.760 0.000 52.300 1.120 ;
  LAYER metal1 ;
  RECT 48.760 0.000 52.300 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 40.080 0.000 43.620 1.120 ;
  LAYER metal3 ;
  RECT 40.080 0.000 43.620 1.120 ;
  LAYER metal2 ;
  RECT 40.080 0.000 43.620 1.120 ;
  LAYER metal1 ;
  RECT 40.080 0.000 43.620 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal3 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal2 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal1 ;
  RECT 27.060 0.000 30.600 1.120 ;
 END
END GND
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 1897.940 125.780 1899.060 129.020 ;
  LAYER metal3 ;
  RECT 1897.940 125.780 1899.060 129.020 ;
  LAYER metal2 ;
  RECT 1897.940 125.780 1899.060 129.020 ;
  LAYER metal1 ;
  RECT 1897.940 125.780 1899.060 129.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1897.940 117.940 1899.060 121.180 ;
  LAYER metal3 ;
  RECT 1897.940 117.940 1899.060 121.180 ;
  LAYER metal2 ;
  RECT 1897.940 117.940 1899.060 121.180 ;
  LAYER metal1 ;
  RECT 1897.940 117.940 1899.060 121.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1897.940 110.100 1899.060 113.340 ;
  LAYER metal3 ;
  RECT 1897.940 110.100 1899.060 113.340 ;
  LAYER metal2 ;
  RECT 1897.940 110.100 1899.060 113.340 ;
  LAYER metal1 ;
  RECT 1897.940 110.100 1899.060 113.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1897.940 102.260 1899.060 105.500 ;
  LAYER metal3 ;
  RECT 1897.940 102.260 1899.060 105.500 ;
  LAYER metal2 ;
  RECT 1897.940 102.260 1899.060 105.500 ;
  LAYER metal1 ;
  RECT 1897.940 102.260 1899.060 105.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1897.940 94.420 1899.060 97.660 ;
  LAYER metal3 ;
  RECT 1897.940 94.420 1899.060 97.660 ;
  LAYER metal2 ;
  RECT 1897.940 94.420 1899.060 97.660 ;
  LAYER metal1 ;
  RECT 1897.940 94.420 1899.060 97.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1897.940 86.580 1899.060 89.820 ;
  LAYER metal3 ;
  RECT 1897.940 86.580 1899.060 89.820 ;
  LAYER metal2 ;
  RECT 1897.940 86.580 1899.060 89.820 ;
  LAYER metal1 ;
  RECT 1897.940 86.580 1899.060 89.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1897.940 47.380 1899.060 50.620 ;
  LAYER metal3 ;
  RECT 1897.940 47.380 1899.060 50.620 ;
  LAYER metal2 ;
  RECT 1897.940 47.380 1899.060 50.620 ;
  LAYER metal1 ;
  RECT 1897.940 47.380 1899.060 50.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1897.940 39.540 1899.060 42.780 ;
  LAYER metal3 ;
  RECT 1897.940 39.540 1899.060 42.780 ;
  LAYER metal2 ;
  RECT 1897.940 39.540 1899.060 42.780 ;
  LAYER metal1 ;
  RECT 1897.940 39.540 1899.060 42.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1897.940 31.700 1899.060 34.940 ;
  LAYER metal3 ;
  RECT 1897.940 31.700 1899.060 34.940 ;
  LAYER metal2 ;
  RECT 1897.940 31.700 1899.060 34.940 ;
  LAYER metal1 ;
  RECT 1897.940 31.700 1899.060 34.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1897.940 23.860 1899.060 27.100 ;
  LAYER metal3 ;
  RECT 1897.940 23.860 1899.060 27.100 ;
  LAYER metal2 ;
  RECT 1897.940 23.860 1899.060 27.100 ;
  LAYER metal1 ;
  RECT 1897.940 23.860 1899.060 27.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1897.940 16.020 1899.060 19.260 ;
  LAYER metal3 ;
  RECT 1897.940 16.020 1899.060 19.260 ;
  LAYER metal2 ;
  RECT 1897.940 16.020 1899.060 19.260 ;
  LAYER metal1 ;
  RECT 1897.940 16.020 1899.060 19.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1897.940 8.180 1899.060 11.420 ;
  LAYER metal3 ;
  RECT 1897.940 8.180 1899.060 11.420 ;
  LAYER metal2 ;
  RECT 1897.940 8.180 1899.060 11.420 ;
  LAYER metal1 ;
  RECT 1897.940 8.180 1899.060 11.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal3 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal2 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal1 ;
  RECT 0.000 125.780 1.120 129.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal3 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal2 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal1 ;
  RECT 0.000 117.940 1.120 121.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal3 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal2 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal1 ;
  RECT 0.000 110.100 1.120 113.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal3 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal2 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal1 ;
  RECT 0.000 102.260 1.120 105.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal3 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal2 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal1 ;
  RECT 0.000 94.420 1.120 97.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal3 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal2 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal1 ;
  RECT 0.000 86.580 1.120 89.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal3 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal2 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal1 ;
  RECT 0.000 47.380 1.120 50.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal3 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal2 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal1 ;
  RECT 0.000 39.540 1.120 42.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal3 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal2 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal1 ;
  RECT 0.000 31.700 1.120 34.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal3 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal2 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal1 ;
  RECT 0.000 23.860 1.120 27.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal3 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal2 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal1 ;
  RECT 0.000 16.020 1.120 19.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal3 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal2 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal1 ;
  RECT 0.000 8.180 1.120 11.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1874.040 165.760 1877.580 166.880 ;
  LAYER metal3 ;
  RECT 1874.040 165.760 1877.580 166.880 ;
  LAYER metal2 ;
  RECT 1874.040 165.760 1877.580 166.880 ;
  LAYER metal1 ;
  RECT 1874.040 165.760 1877.580 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1865.360 165.760 1868.900 166.880 ;
  LAYER metal3 ;
  RECT 1865.360 165.760 1868.900 166.880 ;
  LAYER metal2 ;
  RECT 1865.360 165.760 1868.900 166.880 ;
  LAYER metal1 ;
  RECT 1865.360 165.760 1868.900 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1856.680 165.760 1860.220 166.880 ;
  LAYER metal3 ;
  RECT 1856.680 165.760 1860.220 166.880 ;
  LAYER metal2 ;
  RECT 1856.680 165.760 1860.220 166.880 ;
  LAYER metal1 ;
  RECT 1856.680 165.760 1860.220 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1848.000 165.760 1851.540 166.880 ;
  LAYER metal3 ;
  RECT 1848.000 165.760 1851.540 166.880 ;
  LAYER metal2 ;
  RECT 1848.000 165.760 1851.540 166.880 ;
  LAYER metal1 ;
  RECT 1848.000 165.760 1851.540 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1839.320 165.760 1842.860 166.880 ;
  LAYER metal3 ;
  RECT 1839.320 165.760 1842.860 166.880 ;
  LAYER metal2 ;
  RECT 1839.320 165.760 1842.860 166.880 ;
  LAYER metal1 ;
  RECT 1839.320 165.760 1842.860 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1830.640 165.760 1834.180 166.880 ;
  LAYER metal3 ;
  RECT 1830.640 165.760 1834.180 166.880 ;
  LAYER metal2 ;
  RECT 1830.640 165.760 1834.180 166.880 ;
  LAYER metal1 ;
  RECT 1830.640 165.760 1834.180 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1787.240 165.760 1790.780 166.880 ;
  LAYER metal3 ;
  RECT 1787.240 165.760 1790.780 166.880 ;
  LAYER metal2 ;
  RECT 1787.240 165.760 1790.780 166.880 ;
  LAYER metal1 ;
  RECT 1787.240 165.760 1790.780 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1778.560 165.760 1782.100 166.880 ;
  LAYER metal3 ;
  RECT 1778.560 165.760 1782.100 166.880 ;
  LAYER metal2 ;
  RECT 1778.560 165.760 1782.100 166.880 ;
  LAYER metal1 ;
  RECT 1778.560 165.760 1782.100 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1769.880 165.760 1773.420 166.880 ;
  LAYER metal3 ;
  RECT 1769.880 165.760 1773.420 166.880 ;
  LAYER metal2 ;
  RECT 1769.880 165.760 1773.420 166.880 ;
  LAYER metal1 ;
  RECT 1769.880 165.760 1773.420 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1761.200 165.760 1764.740 166.880 ;
  LAYER metal3 ;
  RECT 1761.200 165.760 1764.740 166.880 ;
  LAYER metal2 ;
  RECT 1761.200 165.760 1764.740 166.880 ;
  LAYER metal1 ;
  RECT 1761.200 165.760 1764.740 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1752.520 165.760 1756.060 166.880 ;
  LAYER metal3 ;
  RECT 1752.520 165.760 1756.060 166.880 ;
  LAYER metal2 ;
  RECT 1752.520 165.760 1756.060 166.880 ;
  LAYER metal1 ;
  RECT 1752.520 165.760 1756.060 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1743.840 165.760 1747.380 166.880 ;
  LAYER metal3 ;
  RECT 1743.840 165.760 1747.380 166.880 ;
  LAYER metal2 ;
  RECT 1743.840 165.760 1747.380 166.880 ;
  LAYER metal1 ;
  RECT 1743.840 165.760 1747.380 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1700.440 165.760 1703.980 166.880 ;
  LAYER metal3 ;
  RECT 1700.440 165.760 1703.980 166.880 ;
  LAYER metal2 ;
  RECT 1700.440 165.760 1703.980 166.880 ;
  LAYER metal1 ;
  RECT 1700.440 165.760 1703.980 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1691.760 165.760 1695.300 166.880 ;
  LAYER metal3 ;
  RECT 1691.760 165.760 1695.300 166.880 ;
  LAYER metal2 ;
  RECT 1691.760 165.760 1695.300 166.880 ;
  LAYER metal1 ;
  RECT 1691.760 165.760 1695.300 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1683.080 165.760 1686.620 166.880 ;
  LAYER metal3 ;
  RECT 1683.080 165.760 1686.620 166.880 ;
  LAYER metal2 ;
  RECT 1683.080 165.760 1686.620 166.880 ;
  LAYER metal1 ;
  RECT 1683.080 165.760 1686.620 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1674.400 165.760 1677.940 166.880 ;
  LAYER metal3 ;
  RECT 1674.400 165.760 1677.940 166.880 ;
  LAYER metal2 ;
  RECT 1674.400 165.760 1677.940 166.880 ;
  LAYER metal1 ;
  RECT 1674.400 165.760 1677.940 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1665.720 165.760 1669.260 166.880 ;
  LAYER metal3 ;
  RECT 1665.720 165.760 1669.260 166.880 ;
  LAYER metal2 ;
  RECT 1665.720 165.760 1669.260 166.880 ;
  LAYER metal1 ;
  RECT 1665.720 165.760 1669.260 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1657.040 165.760 1660.580 166.880 ;
  LAYER metal3 ;
  RECT 1657.040 165.760 1660.580 166.880 ;
  LAYER metal2 ;
  RECT 1657.040 165.760 1660.580 166.880 ;
  LAYER metal1 ;
  RECT 1657.040 165.760 1660.580 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1613.640 165.760 1617.180 166.880 ;
  LAYER metal3 ;
  RECT 1613.640 165.760 1617.180 166.880 ;
  LAYER metal2 ;
  RECT 1613.640 165.760 1617.180 166.880 ;
  LAYER metal1 ;
  RECT 1613.640 165.760 1617.180 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1604.960 165.760 1608.500 166.880 ;
  LAYER metal3 ;
  RECT 1604.960 165.760 1608.500 166.880 ;
  LAYER metal2 ;
  RECT 1604.960 165.760 1608.500 166.880 ;
  LAYER metal1 ;
  RECT 1604.960 165.760 1608.500 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1596.280 165.760 1599.820 166.880 ;
  LAYER metal3 ;
  RECT 1596.280 165.760 1599.820 166.880 ;
  LAYER metal2 ;
  RECT 1596.280 165.760 1599.820 166.880 ;
  LAYER metal1 ;
  RECT 1596.280 165.760 1599.820 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1587.600 165.760 1591.140 166.880 ;
  LAYER metal3 ;
  RECT 1587.600 165.760 1591.140 166.880 ;
  LAYER metal2 ;
  RECT 1587.600 165.760 1591.140 166.880 ;
  LAYER metal1 ;
  RECT 1587.600 165.760 1591.140 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1578.920 165.760 1582.460 166.880 ;
  LAYER metal3 ;
  RECT 1578.920 165.760 1582.460 166.880 ;
  LAYER metal2 ;
  RECT 1578.920 165.760 1582.460 166.880 ;
  LAYER metal1 ;
  RECT 1578.920 165.760 1582.460 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1570.240 165.760 1573.780 166.880 ;
  LAYER metal3 ;
  RECT 1570.240 165.760 1573.780 166.880 ;
  LAYER metal2 ;
  RECT 1570.240 165.760 1573.780 166.880 ;
  LAYER metal1 ;
  RECT 1570.240 165.760 1573.780 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1526.840 165.760 1530.380 166.880 ;
  LAYER metal3 ;
  RECT 1526.840 165.760 1530.380 166.880 ;
  LAYER metal2 ;
  RECT 1526.840 165.760 1530.380 166.880 ;
  LAYER metal1 ;
  RECT 1526.840 165.760 1530.380 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1518.160 165.760 1521.700 166.880 ;
  LAYER metal3 ;
  RECT 1518.160 165.760 1521.700 166.880 ;
  LAYER metal2 ;
  RECT 1518.160 165.760 1521.700 166.880 ;
  LAYER metal1 ;
  RECT 1518.160 165.760 1521.700 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1509.480 165.760 1513.020 166.880 ;
  LAYER metal3 ;
  RECT 1509.480 165.760 1513.020 166.880 ;
  LAYER metal2 ;
  RECT 1509.480 165.760 1513.020 166.880 ;
  LAYER metal1 ;
  RECT 1509.480 165.760 1513.020 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1500.800 165.760 1504.340 166.880 ;
  LAYER metal3 ;
  RECT 1500.800 165.760 1504.340 166.880 ;
  LAYER metal2 ;
  RECT 1500.800 165.760 1504.340 166.880 ;
  LAYER metal1 ;
  RECT 1500.800 165.760 1504.340 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1492.120 165.760 1495.660 166.880 ;
  LAYER metal3 ;
  RECT 1492.120 165.760 1495.660 166.880 ;
  LAYER metal2 ;
  RECT 1492.120 165.760 1495.660 166.880 ;
  LAYER metal1 ;
  RECT 1492.120 165.760 1495.660 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1483.440 165.760 1486.980 166.880 ;
  LAYER metal3 ;
  RECT 1483.440 165.760 1486.980 166.880 ;
  LAYER metal2 ;
  RECT 1483.440 165.760 1486.980 166.880 ;
  LAYER metal1 ;
  RECT 1483.440 165.760 1486.980 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1440.040 165.760 1443.580 166.880 ;
  LAYER metal3 ;
  RECT 1440.040 165.760 1443.580 166.880 ;
  LAYER metal2 ;
  RECT 1440.040 165.760 1443.580 166.880 ;
  LAYER metal1 ;
  RECT 1440.040 165.760 1443.580 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1431.360 165.760 1434.900 166.880 ;
  LAYER metal3 ;
  RECT 1431.360 165.760 1434.900 166.880 ;
  LAYER metal2 ;
  RECT 1431.360 165.760 1434.900 166.880 ;
  LAYER metal1 ;
  RECT 1431.360 165.760 1434.900 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1422.680 165.760 1426.220 166.880 ;
  LAYER metal3 ;
  RECT 1422.680 165.760 1426.220 166.880 ;
  LAYER metal2 ;
  RECT 1422.680 165.760 1426.220 166.880 ;
  LAYER metal1 ;
  RECT 1422.680 165.760 1426.220 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1414.000 165.760 1417.540 166.880 ;
  LAYER metal3 ;
  RECT 1414.000 165.760 1417.540 166.880 ;
  LAYER metal2 ;
  RECT 1414.000 165.760 1417.540 166.880 ;
  LAYER metal1 ;
  RECT 1414.000 165.760 1417.540 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1405.320 165.760 1408.860 166.880 ;
  LAYER metal3 ;
  RECT 1405.320 165.760 1408.860 166.880 ;
  LAYER metal2 ;
  RECT 1405.320 165.760 1408.860 166.880 ;
  LAYER metal1 ;
  RECT 1405.320 165.760 1408.860 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1396.640 165.760 1400.180 166.880 ;
  LAYER metal3 ;
  RECT 1396.640 165.760 1400.180 166.880 ;
  LAYER metal2 ;
  RECT 1396.640 165.760 1400.180 166.880 ;
  LAYER metal1 ;
  RECT 1396.640 165.760 1400.180 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1353.240 165.760 1356.780 166.880 ;
  LAYER metal3 ;
  RECT 1353.240 165.760 1356.780 166.880 ;
  LAYER metal2 ;
  RECT 1353.240 165.760 1356.780 166.880 ;
  LAYER metal1 ;
  RECT 1353.240 165.760 1356.780 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1344.560 165.760 1348.100 166.880 ;
  LAYER metal3 ;
  RECT 1344.560 165.760 1348.100 166.880 ;
  LAYER metal2 ;
  RECT 1344.560 165.760 1348.100 166.880 ;
  LAYER metal1 ;
  RECT 1344.560 165.760 1348.100 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1335.880 165.760 1339.420 166.880 ;
  LAYER metal3 ;
  RECT 1335.880 165.760 1339.420 166.880 ;
  LAYER metal2 ;
  RECT 1335.880 165.760 1339.420 166.880 ;
  LAYER metal1 ;
  RECT 1335.880 165.760 1339.420 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1327.200 165.760 1330.740 166.880 ;
  LAYER metal3 ;
  RECT 1327.200 165.760 1330.740 166.880 ;
  LAYER metal2 ;
  RECT 1327.200 165.760 1330.740 166.880 ;
  LAYER metal1 ;
  RECT 1327.200 165.760 1330.740 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1318.520 165.760 1322.060 166.880 ;
  LAYER metal3 ;
  RECT 1318.520 165.760 1322.060 166.880 ;
  LAYER metal2 ;
  RECT 1318.520 165.760 1322.060 166.880 ;
  LAYER metal1 ;
  RECT 1318.520 165.760 1322.060 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1309.840 165.760 1313.380 166.880 ;
  LAYER metal3 ;
  RECT 1309.840 165.760 1313.380 166.880 ;
  LAYER metal2 ;
  RECT 1309.840 165.760 1313.380 166.880 ;
  LAYER metal1 ;
  RECT 1309.840 165.760 1313.380 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1266.440 165.760 1269.980 166.880 ;
  LAYER metal3 ;
  RECT 1266.440 165.760 1269.980 166.880 ;
  LAYER metal2 ;
  RECT 1266.440 165.760 1269.980 166.880 ;
  LAYER metal1 ;
  RECT 1266.440 165.760 1269.980 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1257.760 165.760 1261.300 166.880 ;
  LAYER metal3 ;
  RECT 1257.760 165.760 1261.300 166.880 ;
  LAYER metal2 ;
  RECT 1257.760 165.760 1261.300 166.880 ;
  LAYER metal1 ;
  RECT 1257.760 165.760 1261.300 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1249.080 165.760 1252.620 166.880 ;
  LAYER metal3 ;
  RECT 1249.080 165.760 1252.620 166.880 ;
  LAYER metal2 ;
  RECT 1249.080 165.760 1252.620 166.880 ;
  LAYER metal1 ;
  RECT 1249.080 165.760 1252.620 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1240.400 165.760 1243.940 166.880 ;
  LAYER metal3 ;
  RECT 1240.400 165.760 1243.940 166.880 ;
  LAYER metal2 ;
  RECT 1240.400 165.760 1243.940 166.880 ;
  LAYER metal1 ;
  RECT 1240.400 165.760 1243.940 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1231.720 165.760 1235.260 166.880 ;
  LAYER metal3 ;
  RECT 1231.720 165.760 1235.260 166.880 ;
  LAYER metal2 ;
  RECT 1231.720 165.760 1235.260 166.880 ;
  LAYER metal1 ;
  RECT 1231.720 165.760 1235.260 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1223.040 165.760 1226.580 166.880 ;
  LAYER metal3 ;
  RECT 1223.040 165.760 1226.580 166.880 ;
  LAYER metal2 ;
  RECT 1223.040 165.760 1226.580 166.880 ;
  LAYER metal1 ;
  RECT 1223.040 165.760 1226.580 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1179.640 165.760 1183.180 166.880 ;
  LAYER metal3 ;
  RECT 1179.640 165.760 1183.180 166.880 ;
  LAYER metal2 ;
  RECT 1179.640 165.760 1183.180 166.880 ;
  LAYER metal1 ;
  RECT 1179.640 165.760 1183.180 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1170.960 165.760 1174.500 166.880 ;
  LAYER metal3 ;
  RECT 1170.960 165.760 1174.500 166.880 ;
  LAYER metal2 ;
  RECT 1170.960 165.760 1174.500 166.880 ;
  LAYER metal1 ;
  RECT 1170.960 165.760 1174.500 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1162.280 165.760 1165.820 166.880 ;
  LAYER metal3 ;
  RECT 1162.280 165.760 1165.820 166.880 ;
  LAYER metal2 ;
  RECT 1162.280 165.760 1165.820 166.880 ;
  LAYER metal1 ;
  RECT 1162.280 165.760 1165.820 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1153.600 165.760 1157.140 166.880 ;
  LAYER metal3 ;
  RECT 1153.600 165.760 1157.140 166.880 ;
  LAYER metal2 ;
  RECT 1153.600 165.760 1157.140 166.880 ;
  LAYER metal1 ;
  RECT 1153.600 165.760 1157.140 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1144.920 165.760 1148.460 166.880 ;
  LAYER metal3 ;
  RECT 1144.920 165.760 1148.460 166.880 ;
  LAYER metal2 ;
  RECT 1144.920 165.760 1148.460 166.880 ;
  LAYER metal1 ;
  RECT 1144.920 165.760 1148.460 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1136.240 165.760 1139.780 166.880 ;
  LAYER metal3 ;
  RECT 1136.240 165.760 1139.780 166.880 ;
  LAYER metal2 ;
  RECT 1136.240 165.760 1139.780 166.880 ;
  LAYER metal1 ;
  RECT 1136.240 165.760 1139.780 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1092.840 165.760 1096.380 166.880 ;
  LAYER metal3 ;
  RECT 1092.840 165.760 1096.380 166.880 ;
  LAYER metal2 ;
  RECT 1092.840 165.760 1096.380 166.880 ;
  LAYER metal1 ;
  RECT 1092.840 165.760 1096.380 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1084.160 165.760 1087.700 166.880 ;
  LAYER metal3 ;
  RECT 1084.160 165.760 1087.700 166.880 ;
  LAYER metal2 ;
  RECT 1084.160 165.760 1087.700 166.880 ;
  LAYER metal1 ;
  RECT 1084.160 165.760 1087.700 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1075.480 165.760 1079.020 166.880 ;
  LAYER metal3 ;
  RECT 1075.480 165.760 1079.020 166.880 ;
  LAYER metal2 ;
  RECT 1075.480 165.760 1079.020 166.880 ;
  LAYER metal1 ;
  RECT 1075.480 165.760 1079.020 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1066.800 165.760 1070.340 166.880 ;
  LAYER metal3 ;
  RECT 1066.800 165.760 1070.340 166.880 ;
  LAYER metal2 ;
  RECT 1066.800 165.760 1070.340 166.880 ;
  LAYER metal1 ;
  RECT 1066.800 165.760 1070.340 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1058.120 165.760 1061.660 166.880 ;
  LAYER metal3 ;
  RECT 1058.120 165.760 1061.660 166.880 ;
  LAYER metal2 ;
  RECT 1058.120 165.760 1061.660 166.880 ;
  LAYER metal1 ;
  RECT 1058.120 165.760 1061.660 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1049.440 165.760 1052.980 166.880 ;
  LAYER metal3 ;
  RECT 1049.440 165.760 1052.980 166.880 ;
  LAYER metal2 ;
  RECT 1049.440 165.760 1052.980 166.880 ;
  LAYER metal1 ;
  RECT 1049.440 165.760 1052.980 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1006.040 165.760 1009.580 166.880 ;
  LAYER metal3 ;
  RECT 1006.040 165.760 1009.580 166.880 ;
  LAYER metal2 ;
  RECT 1006.040 165.760 1009.580 166.880 ;
  LAYER metal1 ;
  RECT 1006.040 165.760 1009.580 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 997.360 165.760 1000.900 166.880 ;
  LAYER metal3 ;
  RECT 997.360 165.760 1000.900 166.880 ;
  LAYER metal2 ;
  RECT 997.360 165.760 1000.900 166.880 ;
  LAYER metal1 ;
  RECT 997.360 165.760 1000.900 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 988.680 165.760 992.220 166.880 ;
  LAYER metal3 ;
  RECT 988.680 165.760 992.220 166.880 ;
  LAYER metal2 ;
  RECT 988.680 165.760 992.220 166.880 ;
  LAYER metal1 ;
  RECT 988.680 165.760 992.220 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 980.000 165.760 983.540 166.880 ;
  LAYER metal3 ;
  RECT 980.000 165.760 983.540 166.880 ;
  LAYER metal2 ;
  RECT 980.000 165.760 983.540 166.880 ;
  LAYER metal1 ;
  RECT 980.000 165.760 983.540 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 971.320 165.760 974.860 166.880 ;
  LAYER metal3 ;
  RECT 971.320 165.760 974.860 166.880 ;
  LAYER metal2 ;
  RECT 971.320 165.760 974.860 166.880 ;
  LAYER metal1 ;
  RECT 971.320 165.760 974.860 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 962.640 165.760 966.180 166.880 ;
  LAYER metal3 ;
  RECT 962.640 165.760 966.180 166.880 ;
  LAYER metal2 ;
  RECT 962.640 165.760 966.180 166.880 ;
  LAYER metal1 ;
  RECT 962.640 165.760 966.180 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 919.240 165.760 922.780 166.880 ;
  LAYER metal3 ;
  RECT 919.240 165.760 922.780 166.880 ;
  LAYER metal2 ;
  RECT 919.240 165.760 922.780 166.880 ;
  LAYER metal1 ;
  RECT 919.240 165.760 922.780 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 910.560 165.760 914.100 166.880 ;
  LAYER metal3 ;
  RECT 910.560 165.760 914.100 166.880 ;
  LAYER metal2 ;
  RECT 910.560 165.760 914.100 166.880 ;
  LAYER metal1 ;
  RECT 910.560 165.760 914.100 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 901.880 165.760 905.420 166.880 ;
  LAYER metal3 ;
  RECT 901.880 165.760 905.420 166.880 ;
  LAYER metal2 ;
  RECT 901.880 165.760 905.420 166.880 ;
  LAYER metal1 ;
  RECT 901.880 165.760 905.420 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 893.200 165.760 896.740 166.880 ;
  LAYER metal3 ;
  RECT 893.200 165.760 896.740 166.880 ;
  LAYER metal2 ;
  RECT 893.200 165.760 896.740 166.880 ;
  LAYER metal1 ;
  RECT 893.200 165.760 896.740 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 884.520 165.760 888.060 166.880 ;
  LAYER metal3 ;
  RECT 884.520 165.760 888.060 166.880 ;
  LAYER metal2 ;
  RECT 884.520 165.760 888.060 166.880 ;
  LAYER metal1 ;
  RECT 884.520 165.760 888.060 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 875.840 165.760 879.380 166.880 ;
  LAYER metal3 ;
  RECT 875.840 165.760 879.380 166.880 ;
  LAYER metal2 ;
  RECT 875.840 165.760 879.380 166.880 ;
  LAYER metal1 ;
  RECT 875.840 165.760 879.380 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 832.440 165.760 835.980 166.880 ;
  LAYER metal3 ;
  RECT 832.440 165.760 835.980 166.880 ;
  LAYER metal2 ;
  RECT 832.440 165.760 835.980 166.880 ;
  LAYER metal1 ;
  RECT 832.440 165.760 835.980 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 823.760 165.760 827.300 166.880 ;
  LAYER metal3 ;
  RECT 823.760 165.760 827.300 166.880 ;
  LAYER metal2 ;
  RECT 823.760 165.760 827.300 166.880 ;
  LAYER metal1 ;
  RECT 823.760 165.760 827.300 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 815.080 165.760 818.620 166.880 ;
  LAYER metal3 ;
  RECT 815.080 165.760 818.620 166.880 ;
  LAYER metal2 ;
  RECT 815.080 165.760 818.620 166.880 ;
  LAYER metal1 ;
  RECT 815.080 165.760 818.620 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 806.400 165.760 809.940 166.880 ;
  LAYER metal3 ;
  RECT 806.400 165.760 809.940 166.880 ;
  LAYER metal2 ;
  RECT 806.400 165.760 809.940 166.880 ;
  LAYER metal1 ;
  RECT 806.400 165.760 809.940 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 797.720 165.760 801.260 166.880 ;
  LAYER metal3 ;
  RECT 797.720 165.760 801.260 166.880 ;
  LAYER metal2 ;
  RECT 797.720 165.760 801.260 166.880 ;
  LAYER metal1 ;
  RECT 797.720 165.760 801.260 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 789.040 165.760 792.580 166.880 ;
  LAYER metal3 ;
  RECT 789.040 165.760 792.580 166.880 ;
  LAYER metal2 ;
  RECT 789.040 165.760 792.580 166.880 ;
  LAYER metal1 ;
  RECT 789.040 165.760 792.580 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 745.640 165.760 749.180 166.880 ;
  LAYER metal3 ;
  RECT 745.640 165.760 749.180 166.880 ;
  LAYER metal2 ;
  RECT 745.640 165.760 749.180 166.880 ;
  LAYER metal1 ;
  RECT 745.640 165.760 749.180 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 736.960 165.760 740.500 166.880 ;
  LAYER metal3 ;
  RECT 736.960 165.760 740.500 166.880 ;
  LAYER metal2 ;
  RECT 736.960 165.760 740.500 166.880 ;
  LAYER metal1 ;
  RECT 736.960 165.760 740.500 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 728.280 165.760 731.820 166.880 ;
  LAYER metal3 ;
  RECT 728.280 165.760 731.820 166.880 ;
  LAYER metal2 ;
  RECT 728.280 165.760 731.820 166.880 ;
  LAYER metal1 ;
  RECT 728.280 165.760 731.820 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 719.600 165.760 723.140 166.880 ;
  LAYER metal3 ;
  RECT 719.600 165.760 723.140 166.880 ;
  LAYER metal2 ;
  RECT 719.600 165.760 723.140 166.880 ;
  LAYER metal1 ;
  RECT 719.600 165.760 723.140 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 710.920 165.760 714.460 166.880 ;
  LAYER metal3 ;
  RECT 710.920 165.760 714.460 166.880 ;
  LAYER metal2 ;
  RECT 710.920 165.760 714.460 166.880 ;
  LAYER metal1 ;
  RECT 710.920 165.760 714.460 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 702.240 165.760 705.780 166.880 ;
  LAYER metal3 ;
  RECT 702.240 165.760 705.780 166.880 ;
  LAYER metal2 ;
  RECT 702.240 165.760 705.780 166.880 ;
  LAYER metal1 ;
  RECT 702.240 165.760 705.780 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 658.840 165.760 662.380 166.880 ;
  LAYER metal3 ;
  RECT 658.840 165.760 662.380 166.880 ;
  LAYER metal2 ;
  RECT 658.840 165.760 662.380 166.880 ;
  LAYER metal1 ;
  RECT 658.840 165.760 662.380 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 650.160 165.760 653.700 166.880 ;
  LAYER metal3 ;
  RECT 650.160 165.760 653.700 166.880 ;
  LAYER metal2 ;
  RECT 650.160 165.760 653.700 166.880 ;
  LAYER metal1 ;
  RECT 650.160 165.760 653.700 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 641.480 165.760 645.020 166.880 ;
  LAYER metal3 ;
  RECT 641.480 165.760 645.020 166.880 ;
  LAYER metal2 ;
  RECT 641.480 165.760 645.020 166.880 ;
  LAYER metal1 ;
  RECT 641.480 165.760 645.020 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 632.800 165.760 636.340 166.880 ;
  LAYER metal3 ;
  RECT 632.800 165.760 636.340 166.880 ;
  LAYER metal2 ;
  RECT 632.800 165.760 636.340 166.880 ;
  LAYER metal1 ;
  RECT 632.800 165.760 636.340 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 624.120 165.760 627.660 166.880 ;
  LAYER metal3 ;
  RECT 624.120 165.760 627.660 166.880 ;
  LAYER metal2 ;
  RECT 624.120 165.760 627.660 166.880 ;
  LAYER metal1 ;
  RECT 624.120 165.760 627.660 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 615.440 165.760 618.980 166.880 ;
  LAYER metal3 ;
  RECT 615.440 165.760 618.980 166.880 ;
  LAYER metal2 ;
  RECT 615.440 165.760 618.980 166.880 ;
  LAYER metal1 ;
  RECT 615.440 165.760 618.980 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 572.040 165.760 575.580 166.880 ;
  LAYER metal3 ;
  RECT 572.040 165.760 575.580 166.880 ;
  LAYER metal2 ;
  RECT 572.040 165.760 575.580 166.880 ;
  LAYER metal1 ;
  RECT 572.040 165.760 575.580 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 563.360 165.760 566.900 166.880 ;
  LAYER metal3 ;
  RECT 563.360 165.760 566.900 166.880 ;
  LAYER metal2 ;
  RECT 563.360 165.760 566.900 166.880 ;
  LAYER metal1 ;
  RECT 563.360 165.760 566.900 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 554.680 165.760 558.220 166.880 ;
  LAYER metal3 ;
  RECT 554.680 165.760 558.220 166.880 ;
  LAYER metal2 ;
  RECT 554.680 165.760 558.220 166.880 ;
  LAYER metal1 ;
  RECT 554.680 165.760 558.220 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 546.000 165.760 549.540 166.880 ;
  LAYER metal3 ;
  RECT 546.000 165.760 549.540 166.880 ;
  LAYER metal2 ;
  RECT 546.000 165.760 549.540 166.880 ;
  LAYER metal1 ;
  RECT 546.000 165.760 549.540 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 537.320 165.760 540.860 166.880 ;
  LAYER metal3 ;
  RECT 537.320 165.760 540.860 166.880 ;
  LAYER metal2 ;
  RECT 537.320 165.760 540.860 166.880 ;
  LAYER metal1 ;
  RECT 537.320 165.760 540.860 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 528.640 165.760 532.180 166.880 ;
  LAYER metal3 ;
  RECT 528.640 165.760 532.180 166.880 ;
  LAYER metal2 ;
  RECT 528.640 165.760 532.180 166.880 ;
  LAYER metal1 ;
  RECT 528.640 165.760 532.180 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 485.240 165.760 488.780 166.880 ;
  LAYER metal3 ;
  RECT 485.240 165.760 488.780 166.880 ;
  LAYER metal2 ;
  RECT 485.240 165.760 488.780 166.880 ;
  LAYER metal1 ;
  RECT 485.240 165.760 488.780 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 476.560 165.760 480.100 166.880 ;
  LAYER metal3 ;
  RECT 476.560 165.760 480.100 166.880 ;
  LAYER metal2 ;
  RECT 476.560 165.760 480.100 166.880 ;
  LAYER metal1 ;
  RECT 476.560 165.760 480.100 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 467.880 165.760 471.420 166.880 ;
  LAYER metal3 ;
  RECT 467.880 165.760 471.420 166.880 ;
  LAYER metal2 ;
  RECT 467.880 165.760 471.420 166.880 ;
  LAYER metal1 ;
  RECT 467.880 165.760 471.420 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 459.200 165.760 462.740 166.880 ;
  LAYER metal3 ;
  RECT 459.200 165.760 462.740 166.880 ;
  LAYER metal2 ;
  RECT 459.200 165.760 462.740 166.880 ;
  LAYER metal1 ;
  RECT 459.200 165.760 462.740 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 450.520 165.760 454.060 166.880 ;
  LAYER metal3 ;
  RECT 450.520 165.760 454.060 166.880 ;
  LAYER metal2 ;
  RECT 450.520 165.760 454.060 166.880 ;
  LAYER metal1 ;
  RECT 450.520 165.760 454.060 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 441.840 165.760 445.380 166.880 ;
  LAYER metal3 ;
  RECT 441.840 165.760 445.380 166.880 ;
  LAYER metal2 ;
  RECT 441.840 165.760 445.380 166.880 ;
  LAYER metal1 ;
  RECT 441.840 165.760 445.380 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 398.440 165.760 401.980 166.880 ;
  LAYER metal3 ;
  RECT 398.440 165.760 401.980 166.880 ;
  LAYER metal2 ;
  RECT 398.440 165.760 401.980 166.880 ;
  LAYER metal1 ;
  RECT 398.440 165.760 401.980 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 389.760 165.760 393.300 166.880 ;
  LAYER metal3 ;
  RECT 389.760 165.760 393.300 166.880 ;
  LAYER metal2 ;
  RECT 389.760 165.760 393.300 166.880 ;
  LAYER metal1 ;
  RECT 389.760 165.760 393.300 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 381.080 165.760 384.620 166.880 ;
  LAYER metal3 ;
  RECT 381.080 165.760 384.620 166.880 ;
  LAYER metal2 ;
  RECT 381.080 165.760 384.620 166.880 ;
  LAYER metal1 ;
  RECT 381.080 165.760 384.620 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 372.400 165.760 375.940 166.880 ;
  LAYER metal3 ;
  RECT 372.400 165.760 375.940 166.880 ;
  LAYER metal2 ;
  RECT 372.400 165.760 375.940 166.880 ;
  LAYER metal1 ;
  RECT 372.400 165.760 375.940 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 363.720 165.760 367.260 166.880 ;
  LAYER metal3 ;
  RECT 363.720 165.760 367.260 166.880 ;
  LAYER metal2 ;
  RECT 363.720 165.760 367.260 166.880 ;
  LAYER metal1 ;
  RECT 363.720 165.760 367.260 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 355.040 165.760 358.580 166.880 ;
  LAYER metal3 ;
  RECT 355.040 165.760 358.580 166.880 ;
  LAYER metal2 ;
  RECT 355.040 165.760 358.580 166.880 ;
  LAYER metal1 ;
  RECT 355.040 165.760 358.580 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 311.640 165.760 315.180 166.880 ;
  LAYER metal3 ;
  RECT 311.640 165.760 315.180 166.880 ;
  LAYER metal2 ;
  RECT 311.640 165.760 315.180 166.880 ;
  LAYER metal1 ;
  RECT 311.640 165.760 315.180 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 302.960 165.760 306.500 166.880 ;
  LAYER metal3 ;
  RECT 302.960 165.760 306.500 166.880 ;
  LAYER metal2 ;
  RECT 302.960 165.760 306.500 166.880 ;
  LAYER metal1 ;
  RECT 302.960 165.760 306.500 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 294.280 165.760 297.820 166.880 ;
  LAYER metal3 ;
  RECT 294.280 165.760 297.820 166.880 ;
  LAYER metal2 ;
  RECT 294.280 165.760 297.820 166.880 ;
  LAYER metal1 ;
  RECT 294.280 165.760 297.820 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 285.600 165.760 289.140 166.880 ;
  LAYER metal3 ;
  RECT 285.600 165.760 289.140 166.880 ;
  LAYER metal2 ;
  RECT 285.600 165.760 289.140 166.880 ;
  LAYER metal1 ;
  RECT 285.600 165.760 289.140 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 276.920 165.760 280.460 166.880 ;
  LAYER metal3 ;
  RECT 276.920 165.760 280.460 166.880 ;
  LAYER metal2 ;
  RECT 276.920 165.760 280.460 166.880 ;
  LAYER metal1 ;
  RECT 276.920 165.760 280.460 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 268.240 165.760 271.780 166.880 ;
  LAYER metal3 ;
  RECT 268.240 165.760 271.780 166.880 ;
  LAYER metal2 ;
  RECT 268.240 165.760 271.780 166.880 ;
  LAYER metal1 ;
  RECT 268.240 165.760 271.780 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 224.840 165.760 228.380 166.880 ;
  LAYER metal3 ;
  RECT 224.840 165.760 228.380 166.880 ;
  LAYER metal2 ;
  RECT 224.840 165.760 228.380 166.880 ;
  LAYER metal1 ;
  RECT 224.840 165.760 228.380 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 216.160 165.760 219.700 166.880 ;
  LAYER metal3 ;
  RECT 216.160 165.760 219.700 166.880 ;
  LAYER metal2 ;
  RECT 216.160 165.760 219.700 166.880 ;
  LAYER metal1 ;
  RECT 216.160 165.760 219.700 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 207.480 165.760 211.020 166.880 ;
  LAYER metal3 ;
  RECT 207.480 165.760 211.020 166.880 ;
  LAYER metal2 ;
  RECT 207.480 165.760 211.020 166.880 ;
  LAYER metal1 ;
  RECT 207.480 165.760 211.020 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 198.800 165.760 202.340 166.880 ;
  LAYER metal3 ;
  RECT 198.800 165.760 202.340 166.880 ;
  LAYER metal2 ;
  RECT 198.800 165.760 202.340 166.880 ;
  LAYER metal1 ;
  RECT 198.800 165.760 202.340 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 190.120 165.760 193.660 166.880 ;
  LAYER metal3 ;
  RECT 190.120 165.760 193.660 166.880 ;
  LAYER metal2 ;
  RECT 190.120 165.760 193.660 166.880 ;
  LAYER metal1 ;
  RECT 190.120 165.760 193.660 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 181.440 165.760 184.980 166.880 ;
  LAYER metal3 ;
  RECT 181.440 165.760 184.980 166.880 ;
  LAYER metal2 ;
  RECT 181.440 165.760 184.980 166.880 ;
  LAYER metal1 ;
  RECT 181.440 165.760 184.980 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 138.040 165.760 141.580 166.880 ;
  LAYER metal3 ;
  RECT 138.040 165.760 141.580 166.880 ;
  LAYER metal2 ;
  RECT 138.040 165.760 141.580 166.880 ;
  LAYER metal1 ;
  RECT 138.040 165.760 141.580 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 129.360 165.760 132.900 166.880 ;
  LAYER metal3 ;
  RECT 129.360 165.760 132.900 166.880 ;
  LAYER metal2 ;
  RECT 129.360 165.760 132.900 166.880 ;
  LAYER metal1 ;
  RECT 129.360 165.760 132.900 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 120.680 165.760 124.220 166.880 ;
  LAYER metal3 ;
  RECT 120.680 165.760 124.220 166.880 ;
  LAYER metal2 ;
  RECT 120.680 165.760 124.220 166.880 ;
  LAYER metal1 ;
  RECT 120.680 165.760 124.220 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 112.000 165.760 115.540 166.880 ;
  LAYER metal3 ;
  RECT 112.000 165.760 115.540 166.880 ;
  LAYER metal2 ;
  RECT 112.000 165.760 115.540 166.880 ;
  LAYER metal1 ;
  RECT 112.000 165.760 115.540 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 103.320 165.760 106.860 166.880 ;
  LAYER metal3 ;
  RECT 103.320 165.760 106.860 166.880 ;
  LAYER metal2 ;
  RECT 103.320 165.760 106.860 166.880 ;
  LAYER metal1 ;
  RECT 103.320 165.760 106.860 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 94.640 165.760 98.180 166.880 ;
  LAYER metal3 ;
  RECT 94.640 165.760 98.180 166.880 ;
  LAYER metal2 ;
  RECT 94.640 165.760 98.180 166.880 ;
  LAYER metal1 ;
  RECT 94.640 165.760 98.180 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 51.240 165.760 54.780 166.880 ;
  LAYER metal3 ;
  RECT 51.240 165.760 54.780 166.880 ;
  LAYER metal2 ;
  RECT 51.240 165.760 54.780 166.880 ;
  LAYER metal1 ;
  RECT 51.240 165.760 54.780 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 42.560 165.760 46.100 166.880 ;
  LAYER metal3 ;
  RECT 42.560 165.760 46.100 166.880 ;
  LAYER metal2 ;
  RECT 42.560 165.760 46.100 166.880 ;
  LAYER metal1 ;
  RECT 42.560 165.760 46.100 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 33.880 165.760 37.420 166.880 ;
  LAYER metal3 ;
  RECT 33.880 165.760 37.420 166.880 ;
  LAYER metal2 ;
  RECT 33.880 165.760 37.420 166.880 ;
  LAYER metal1 ;
  RECT 33.880 165.760 37.420 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 25.200 165.760 28.740 166.880 ;
  LAYER metal3 ;
  RECT 25.200 165.760 28.740 166.880 ;
  LAYER metal2 ;
  RECT 25.200 165.760 28.740 166.880 ;
  LAYER metal1 ;
  RECT 25.200 165.760 28.740 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 16.520 165.760 20.060 166.880 ;
  LAYER metal3 ;
  RECT 16.520 165.760 20.060 166.880 ;
  LAYER metal2 ;
  RECT 16.520 165.760 20.060 166.880 ;
  LAYER metal1 ;
  RECT 16.520 165.760 20.060 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 7.840 165.760 11.380 166.880 ;
  LAYER metal3 ;
  RECT 7.840 165.760 11.380 166.880 ;
  LAYER metal2 ;
  RECT 7.840 165.760 11.380 166.880 ;
  LAYER metal1 ;
  RECT 7.840 165.760 11.380 166.880 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1852.960 0.000 1856.500 1.120 ;
  LAYER metal3 ;
  RECT 1852.960 0.000 1856.500 1.120 ;
  LAYER metal2 ;
  RECT 1852.960 0.000 1856.500 1.120 ;
  LAYER metal1 ;
  RECT 1852.960 0.000 1856.500 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1844.280 0.000 1847.820 1.120 ;
  LAYER metal3 ;
  RECT 1844.280 0.000 1847.820 1.120 ;
  LAYER metal2 ;
  RECT 1844.280 0.000 1847.820 1.120 ;
  LAYER metal1 ;
  RECT 1844.280 0.000 1847.820 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1835.600 0.000 1839.140 1.120 ;
  LAYER metal3 ;
  RECT 1835.600 0.000 1839.140 1.120 ;
  LAYER metal2 ;
  RECT 1835.600 0.000 1839.140 1.120 ;
  LAYER metal1 ;
  RECT 1835.600 0.000 1839.140 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1826.920 0.000 1830.460 1.120 ;
  LAYER metal3 ;
  RECT 1826.920 0.000 1830.460 1.120 ;
  LAYER metal2 ;
  RECT 1826.920 0.000 1830.460 1.120 ;
  LAYER metal1 ;
  RECT 1826.920 0.000 1830.460 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1818.240 0.000 1821.780 1.120 ;
  LAYER metal3 ;
  RECT 1818.240 0.000 1821.780 1.120 ;
  LAYER metal2 ;
  RECT 1818.240 0.000 1821.780 1.120 ;
  LAYER metal1 ;
  RECT 1818.240 0.000 1821.780 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1809.560 0.000 1813.100 1.120 ;
  LAYER metal3 ;
  RECT 1809.560 0.000 1813.100 1.120 ;
  LAYER metal2 ;
  RECT 1809.560 0.000 1813.100 1.120 ;
  LAYER metal1 ;
  RECT 1809.560 0.000 1813.100 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1748.800 0.000 1752.340 1.120 ;
  LAYER metal3 ;
  RECT 1748.800 0.000 1752.340 1.120 ;
  LAYER metal2 ;
  RECT 1748.800 0.000 1752.340 1.120 ;
  LAYER metal1 ;
  RECT 1748.800 0.000 1752.340 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1740.120 0.000 1743.660 1.120 ;
  LAYER metal3 ;
  RECT 1740.120 0.000 1743.660 1.120 ;
  LAYER metal2 ;
  RECT 1740.120 0.000 1743.660 1.120 ;
  LAYER metal1 ;
  RECT 1740.120 0.000 1743.660 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1731.440 0.000 1734.980 1.120 ;
  LAYER metal3 ;
  RECT 1731.440 0.000 1734.980 1.120 ;
  LAYER metal2 ;
  RECT 1731.440 0.000 1734.980 1.120 ;
  LAYER metal1 ;
  RECT 1731.440 0.000 1734.980 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1722.760 0.000 1726.300 1.120 ;
  LAYER metal3 ;
  RECT 1722.760 0.000 1726.300 1.120 ;
  LAYER metal2 ;
  RECT 1722.760 0.000 1726.300 1.120 ;
  LAYER metal1 ;
  RECT 1722.760 0.000 1726.300 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1714.080 0.000 1717.620 1.120 ;
  LAYER metal3 ;
  RECT 1714.080 0.000 1717.620 1.120 ;
  LAYER metal2 ;
  RECT 1714.080 0.000 1717.620 1.120 ;
  LAYER metal1 ;
  RECT 1714.080 0.000 1717.620 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1705.400 0.000 1708.940 1.120 ;
  LAYER metal3 ;
  RECT 1705.400 0.000 1708.940 1.120 ;
  LAYER metal2 ;
  RECT 1705.400 0.000 1708.940 1.120 ;
  LAYER metal1 ;
  RECT 1705.400 0.000 1708.940 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1644.640 0.000 1648.180 1.120 ;
  LAYER metal3 ;
  RECT 1644.640 0.000 1648.180 1.120 ;
  LAYER metal2 ;
  RECT 1644.640 0.000 1648.180 1.120 ;
  LAYER metal1 ;
  RECT 1644.640 0.000 1648.180 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1635.960 0.000 1639.500 1.120 ;
  LAYER metal3 ;
  RECT 1635.960 0.000 1639.500 1.120 ;
  LAYER metal2 ;
  RECT 1635.960 0.000 1639.500 1.120 ;
  LAYER metal1 ;
  RECT 1635.960 0.000 1639.500 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1627.280 0.000 1630.820 1.120 ;
  LAYER metal3 ;
  RECT 1627.280 0.000 1630.820 1.120 ;
  LAYER metal2 ;
  RECT 1627.280 0.000 1630.820 1.120 ;
  LAYER metal1 ;
  RECT 1627.280 0.000 1630.820 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1618.600 0.000 1622.140 1.120 ;
  LAYER metal3 ;
  RECT 1618.600 0.000 1622.140 1.120 ;
  LAYER metal2 ;
  RECT 1618.600 0.000 1622.140 1.120 ;
  LAYER metal1 ;
  RECT 1618.600 0.000 1622.140 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1609.920 0.000 1613.460 1.120 ;
  LAYER metal3 ;
  RECT 1609.920 0.000 1613.460 1.120 ;
  LAYER metal2 ;
  RECT 1609.920 0.000 1613.460 1.120 ;
  LAYER metal1 ;
  RECT 1609.920 0.000 1613.460 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1601.240 0.000 1604.780 1.120 ;
  LAYER metal3 ;
  RECT 1601.240 0.000 1604.780 1.120 ;
  LAYER metal2 ;
  RECT 1601.240 0.000 1604.780 1.120 ;
  LAYER metal1 ;
  RECT 1601.240 0.000 1604.780 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1539.860 0.000 1543.400 1.120 ;
  LAYER metal3 ;
  RECT 1539.860 0.000 1543.400 1.120 ;
  LAYER metal2 ;
  RECT 1539.860 0.000 1543.400 1.120 ;
  LAYER metal1 ;
  RECT 1539.860 0.000 1543.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1531.180 0.000 1534.720 1.120 ;
  LAYER metal3 ;
  RECT 1531.180 0.000 1534.720 1.120 ;
  LAYER metal2 ;
  RECT 1531.180 0.000 1534.720 1.120 ;
  LAYER metal1 ;
  RECT 1531.180 0.000 1534.720 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1522.500 0.000 1526.040 1.120 ;
  LAYER metal3 ;
  RECT 1522.500 0.000 1526.040 1.120 ;
  LAYER metal2 ;
  RECT 1522.500 0.000 1526.040 1.120 ;
  LAYER metal1 ;
  RECT 1522.500 0.000 1526.040 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1513.820 0.000 1517.360 1.120 ;
  LAYER metal3 ;
  RECT 1513.820 0.000 1517.360 1.120 ;
  LAYER metal2 ;
  RECT 1513.820 0.000 1517.360 1.120 ;
  LAYER metal1 ;
  RECT 1513.820 0.000 1517.360 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1505.140 0.000 1508.680 1.120 ;
  LAYER metal3 ;
  RECT 1505.140 0.000 1508.680 1.120 ;
  LAYER metal2 ;
  RECT 1505.140 0.000 1508.680 1.120 ;
  LAYER metal1 ;
  RECT 1505.140 0.000 1508.680 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1496.460 0.000 1500.000 1.120 ;
  LAYER metal3 ;
  RECT 1496.460 0.000 1500.000 1.120 ;
  LAYER metal2 ;
  RECT 1496.460 0.000 1500.000 1.120 ;
  LAYER metal1 ;
  RECT 1496.460 0.000 1500.000 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1440.040 0.000 1443.580 1.120 ;
  LAYER metal3 ;
  RECT 1440.040 0.000 1443.580 1.120 ;
  LAYER metal2 ;
  RECT 1440.040 0.000 1443.580 1.120 ;
  LAYER metal1 ;
  RECT 1440.040 0.000 1443.580 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1427.020 0.000 1430.560 1.120 ;
  LAYER metal3 ;
  RECT 1427.020 0.000 1430.560 1.120 ;
  LAYER metal2 ;
  RECT 1427.020 0.000 1430.560 1.120 ;
  LAYER metal1 ;
  RECT 1427.020 0.000 1430.560 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1418.340 0.000 1421.880 1.120 ;
  LAYER metal3 ;
  RECT 1418.340 0.000 1421.880 1.120 ;
  LAYER metal2 ;
  RECT 1418.340 0.000 1421.880 1.120 ;
  LAYER metal1 ;
  RECT 1418.340 0.000 1421.880 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1409.660 0.000 1413.200 1.120 ;
  LAYER metal3 ;
  RECT 1409.660 0.000 1413.200 1.120 ;
  LAYER metal2 ;
  RECT 1409.660 0.000 1413.200 1.120 ;
  LAYER metal1 ;
  RECT 1409.660 0.000 1413.200 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1400.980 0.000 1404.520 1.120 ;
  LAYER metal3 ;
  RECT 1400.980 0.000 1404.520 1.120 ;
  LAYER metal2 ;
  RECT 1400.980 0.000 1404.520 1.120 ;
  LAYER metal1 ;
  RECT 1400.980 0.000 1404.520 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1392.300 0.000 1395.840 1.120 ;
  LAYER metal3 ;
  RECT 1392.300 0.000 1395.840 1.120 ;
  LAYER metal2 ;
  RECT 1392.300 0.000 1395.840 1.120 ;
  LAYER metal1 ;
  RECT 1392.300 0.000 1395.840 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1348.900 0.000 1352.440 1.120 ;
  LAYER metal3 ;
  RECT 1348.900 0.000 1352.440 1.120 ;
  LAYER metal2 ;
  RECT 1348.900 0.000 1352.440 1.120 ;
  LAYER metal1 ;
  RECT 1348.900 0.000 1352.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1327.200 0.000 1330.740 1.120 ;
  LAYER metal3 ;
  RECT 1327.200 0.000 1330.740 1.120 ;
  LAYER metal2 ;
  RECT 1327.200 0.000 1330.740 1.120 ;
  LAYER metal1 ;
  RECT 1327.200 0.000 1330.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1314.180 0.000 1317.720 1.120 ;
  LAYER metal3 ;
  RECT 1314.180 0.000 1317.720 1.120 ;
  LAYER metal2 ;
  RECT 1314.180 0.000 1317.720 1.120 ;
  LAYER metal1 ;
  RECT 1314.180 0.000 1317.720 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1305.500 0.000 1309.040 1.120 ;
  LAYER metal3 ;
  RECT 1305.500 0.000 1309.040 1.120 ;
  LAYER metal2 ;
  RECT 1305.500 0.000 1309.040 1.120 ;
  LAYER metal1 ;
  RECT 1305.500 0.000 1309.040 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1296.820 0.000 1300.360 1.120 ;
  LAYER metal3 ;
  RECT 1296.820 0.000 1300.360 1.120 ;
  LAYER metal2 ;
  RECT 1296.820 0.000 1300.360 1.120 ;
  LAYER metal1 ;
  RECT 1296.820 0.000 1300.360 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1288.140 0.000 1291.680 1.120 ;
  LAYER metal3 ;
  RECT 1288.140 0.000 1291.680 1.120 ;
  LAYER metal2 ;
  RECT 1288.140 0.000 1291.680 1.120 ;
  LAYER metal1 ;
  RECT 1288.140 0.000 1291.680 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1244.740 0.000 1248.280 1.120 ;
  LAYER metal3 ;
  RECT 1244.740 0.000 1248.280 1.120 ;
  LAYER metal2 ;
  RECT 1244.740 0.000 1248.280 1.120 ;
  LAYER metal1 ;
  RECT 1244.740 0.000 1248.280 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1236.060 0.000 1239.600 1.120 ;
  LAYER metal3 ;
  RECT 1236.060 0.000 1239.600 1.120 ;
  LAYER metal2 ;
  RECT 1236.060 0.000 1239.600 1.120 ;
  LAYER metal1 ;
  RECT 1236.060 0.000 1239.600 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1214.360 0.000 1217.900 1.120 ;
  LAYER metal3 ;
  RECT 1214.360 0.000 1217.900 1.120 ;
  LAYER metal2 ;
  RECT 1214.360 0.000 1217.900 1.120 ;
  LAYER metal1 ;
  RECT 1214.360 0.000 1217.900 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1200.720 0.000 1204.260 1.120 ;
  LAYER metal3 ;
  RECT 1200.720 0.000 1204.260 1.120 ;
  LAYER metal2 ;
  RECT 1200.720 0.000 1204.260 1.120 ;
  LAYER metal1 ;
  RECT 1200.720 0.000 1204.260 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1192.040 0.000 1195.580 1.120 ;
  LAYER metal3 ;
  RECT 1192.040 0.000 1195.580 1.120 ;
  LAYER metal2 ;
  RECT 1192.040 0.000 1195.580 1.120 ;
  LAYER metal1 ;
  RECT 1192.040 0.000 1195.580 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1183.360 0.000 1186.900 1.120 ;
  LAYER metal3 ;
  RECT 1183.360 0.000 1186.900 1.120 ;
  LAYER metal2 ;
  RECT 1183.360 0.000 1186.900 1.120 ;
  LAYER metal1 ;
  RECT 1183.360 0.000 1186.900 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1139.960 0.000 1143.500 1.120 ;
  LAYER metal3 ;
  RECT 1139.960 0.000 1143.500 1.120 ;
  LAYER metal2 ;
  RECT 1139.960 0.000 1143.500 1.120 ;
  LAYER metal1 ;
  RECT 1139.960 0.000 1143.500 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1131.280 0.000 1134.820 1.120 ;
  LAYER metal3 ;
  RECT 1131.280 0.000 1134.820 1.120 ;
  LAYER metal2 ;
  RECT 1131.280 0.000 1134.820 1.120 ;
  LAYER metal1 ;
  RECT 1131.280 0.000 1134.820 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1122.600 0.000 1126.140 1.120 ;
  LAYER metal3 ;
  RECT 1122.600 0.000 1126.140 1.120 ;
  LAYER metal2 ;
  RECT 1122.600 0.000 1126.140 1.120 ;
  LAYER metal1 ;
  RECT 1122.600 0.000 1126.140 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1100.900 0.000 1104.440 1.120 ;
  LAYER metal3 ;
  RECT 1100.900 0.000 1104.440 1.120 ;
  LAYER metal2 ;
  RECT 1100.900 0.000 1104.440 1.120 ;
  LAYER metal1 ;
  RECT 1100.900 0.000 1104.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1087.880 0.000 1091.420 1.120 ;
  LAYER metal3 ;
  RECT 1087.880 0.000 1091.420 1.120 ;
  LAYER metal2 ;
  RECT 1087.880 0.000 1091.420 1.120 ;
  LAYER metal1 ;
  RECT 1087.880 0.000 1091.420 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1079.200 0.000 1082.740 1.120 ;
  LAYER metal3 ;
  RECT 1079.200 0.000 1082.740 1.120 ;
  LAYER metal2 ;
  RECT 1079.200 0.000 1082.740 1.120 ;
  LAYER metal1 ;
  RECT 1079.200 0.000 1082.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1035.800 0.000 1039.340 1.120 ;
  LAYER metal3 ;
  RECT 1035.800 0.000 1039.340 1.120 ;
  LAYER metal2 ;
  RECT 1035.800 0.000 1039.340 1.120 ;
  LAYER metal1 ;
  RECT 1035.800 0.000 1039.340 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1027.120 0.000 1030.660 1.120 ;
  LAYER metal3 ;
  RECT 1027.120 0.000 1030.660 1.120 ;
  LAYER metal2 ;
  RECT 1027.120 0.000 1030.660 1.120 ;
  LAYER metal1 ;
  RECT 1027.120 0.000 1030.660 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1018.440 0.000 1021.980 1.120 ;
  LAYER metal3 ;
  RECT 1018.440 0.000 1021.980 1.120 ;
  LAYER metal2 ;
  RECT 1018.440 0.000 1021.980 1.120 ;
  LAYER metal1 ;
  RECT 1018.440 0.000 1021.980 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 1009.760 0.000 1013.300 1.120 ;
  LAYER metal3 ;
  RECT 1009.760 0.000 1013.300 1.120 ;
  LAYER metal2 ;
  RECT 1009.760 0.000 1013.300 1.120 ;
  LAYER metal1 ;
  RECT 1009.760 0.000 1013.300 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 988.060 0.000 991.600 1.120 ;
  LAYER metal3 ;
  RECT 988.060 0.000 991.600 1.120 ;
  LAYER metal2 ;
  RECT 988.060 0.000 991.600 1.120 ;
  LAYER metal1 ;
  RECT 988.060 0.000 991.600 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 956.440 0.000 959.980 1.120 ;
  LAYER metal3 ;
  RECT 956.440 0.000 959.980 1.120 ;
  LAYER metal2 ;
  RECT 956.440 0.000 959.980 1.120 ;
  LAYER metal1 ;
  RECT 956.440 0.000 959.980 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 887.620 0.000 891.160 1.120 ;
  LAYER metal3 ;
  RECT 887.620 0.000 891.160 1.120 ;
  LAYER metal2 ;
  RECT 887.620 0.000 891.160 1.120 ;
  LAYER metal1 ;
  RECT 887.620 0.000 891.160 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 878.940 0.000 882.480 1.120 ;
  LAYER metal3 ;
  RECT 878.940 0.000 882.480 1.120 ;
  LAYER metal2 ;
  RECT 878.940 0.000 882.480 1.120 ;
  LAYER metal1 ;
  RECT 878.940 0.000 882.480 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 870.260 0.000 873.800 1.120 ;
  LAYER metal3 ;
  RECT 870.260 0.000 873.800 1.120 ;
  LAYER metal2 ;
  RECT 870.260 0.000 873.800 1.120 ;
  LAYER metal1 ;
  RECT 870.260 0.000 873.800 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 861.580 0.000 865.120 1.120 ;
  LAYER metal3 ;
  RECT 861.580 0.000 865.120 1.120 ;
  LAYER metal2 ;
  RECT 861.580 0.000 865.120 1.120 ;
  LAYER metal1 ;
  RECT 861.580 0.000 865.120 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 852.900 0.000 856.440 1.120 ;
  LAYER metal3 ;
  RECT 852.900 0.000 856.440 1.120 ;
  LAYER metal2 ;
  RECT 852.900 0.000 856.440 1.120 ;
  LAYER metal1 ;
  RECT 852.900 0.000 856.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 844.220 0.000 847.760 1.120 ;
  LAYER metal3 ;
  RECT 844.220 0.000 847.760 1.120 ;
  LAYER metal2 ;
  RECT 844.220 0.000 847.760 1.120 ;
  LAYER metal1 ;
  RECT 844.220 0.000 847.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 783.460 0.000 787.000 1.120 ;
  LAYER metal3 ;
  RECT 783.460 0.000 787.000 1.120 ;
  LAYER metal2 ;
  RECT 783.460 0.000 787.000 1.120 ;
  LAYER metal1 ;
  RECT 783.460 0.000 787.000 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 774.780 0.000 778.320 1.120 ;
  LAYER metal3 ;
  RECT 774.780 0.000 778.320 1.120 ;
  LAYER metal2 ;
  RECT 774.780 0.000 778.320 1.120 ;
  LAYER metal1 ;
  RECT 774.780 0.000 778.320 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 766.100 0.000 769.640 1.120 ;
  LAYER metal3 ;
  RECT 766.100 0.000 769.640 1.120 ;
  LAYER metal2 ;
  RECT 766.100 0.000 769.640 1.120 ;
  LAYER metal1 ;
  RECT 766.100 0.000 769.640 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 757.420 0.000 760.960 1.120 ;
  LAYER metal3 ;
  RECT 757.420 0.000 760.960 1.120 ;
  LAYER metal2 ;
  RECT 757.420 0.000 760.960 1.120 ;
  LAYER metal1 ;
  RECT 757.420 0.000 760.960 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 748.740 0.000 752.280 1.120 ;
  LAYER metal3 ;
  RECT 748.740 0.000 752.280 1.120 ;
  LAYER metal2 ;
  RECT 748.740 0.000 752.280 1.120 ;
  LAYER metal1 ;
  RECT 748.740 0.000 752.280 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 740.060 0.000 743.600 1.120 ;
  LAYER metal3 ;
  RECT 740.060 0.000 743.600 1.120 ;
  LAYER metal2 ;
  RECT 740.060 0.000 743.600 1.120 ;
  LAYER metal1 ;
  RECT 740.060 0.000 743.600 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 678.680 0.000 682.220 1.120 ;
  LAYER metal3 ;
  RECT 678.680 0.000 682.220 1.120 ;
  LAYER metal2 ;
  RECT 678.680 0.000 682.220 1.120 ;
  LAYER metal1 ;
  RECT 678.680 0.000 682.220 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 670.000 0.000 673.540 1.120 ;
  LAYER metal3 ;
  RECT 670.000 0.000 673.540 1.120 ;
  LAYER metal2 ;
  RECT 670.000 0.000 673.540 1.120 ;
  LAYER metal1 ;
  RECT 670.000 0.000 673.540 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 661.320 0.000 664.860 1.120 ;
  LAYER metal3 ;
  RECT 661.320 0.000 664.860 1.120 ;
  LAYER metal2 ;
  RECT 661.320 0.000 664.860 1.120 ;
  LAYER metal1 ;
  RECT 661.320 0.000 664.860 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 652.640 0.000 656.180 1.120 ;
  LAYER metal3 ;
  RECT 652.640 0.000 656.180 1.120 ;
  LAYER metal2 ;
  RECT 652.640 0.000 656.180 1.120 ;
  LAYER metal1 ;
  RECT 652.640 0.000 656.180 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 643.960 0.000 647.500 1.120 ;
  LAYER metal3 ;
  RECT 643.960 0.000 647.500 1.120 ;
  LAYER metal2 ;
  RECT 643.960 0.000 647.500 1.120 ;
  LAYER metal1 ;
  RECT 643.960 0.000 647.500 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 635.280 0.000 638.820 1.120 ;
  LAYER metal3 ;
  RECT 635.280 0.000 638.820 1.120 ;
  LAYER metal2 ;
  RECT 635.280 0.000 638.820 1.120 ;
  LAYER metal1 ;
  RECT 635.280 0.000 638.820 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 578.860 0.000 582.400 1.120 ;
  LAYER metal3 ;
  RECT 578.860 0.000 582.400 1.120 ;
  LAYER metal2 ;
  RECT 578.860 0.000 582.400 1.120 ;
  LAYER metal1 ;
  RECT 578.860 0.000 582.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER metal3 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER metal2 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER metal1 ;
  RECT 565.840 0.000 569.380 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 557.160 0.000 560.700 1.120 ;
  LAYER metal3 ;
  RECT 557.160 0.000 560.700 1.120 ;
  LAYER metal2 ;
  RECT 557.160 0.000 560.700 1.120 ;
  LAYER metal1 ;
  RECT 557.160 0.000 560.700 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 548.480 0.000 552.020 1.120 ;
  LAYER metal3 ;
  RECT 548.480 0.000 552.020 1.120 ;
  LAYER metal2 ;
  RECT 548.480 0.000 552.020 1.120 ;
  LAYER metal1 ;
  RECT 548.480 0.000 552.020 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 539.800 0.000 543.340 1.120 ;
  LAYER metal3 ;
  RECT 539.800 0.000 543.340 1.120 ;
  LAYER metal2 ;
  RECT 539.800 0.000 543.340 1.120 ;
  LAYER metal1 ;
  RECT 539.800 0.000 543.340 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 531.120 0.000 534.660 1.120 ;
  LAYER metal3 ;
  RECT 531.120 0.000 534.660 1.120 ;
  LAYER metal2 ;
  RECT 531.120 0.000 534.660 1.120 ;
  LAYER metal1 ;
  RECT 531.120 0.000 534.660 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 487.720 0.000 491.260 1.120 ;
  LAYER metal3 ;
  RECT 487.720 0.000 491.260 1.120 ;
  LAYER metal2 ;
  RECT 487.720 0.000 491.260 1.120 ;
  LAYER metal1 ;
  RECT 487.720 0.000 491.260 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 466.020 0.000 469.560 1.120 ;
  LAYER metal3 ;
  RECT 466.020 0.000 469.560 1.120 ;
  LAYER metal2 ;
  RECT 466.020 0.000 469.560 1.120 ;
  LAYER metal1 ;
  RECT 466.020 0.000 469.560 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 453.000 0.000 456.540 1.120 ;
  LAYER metal3 ;
  RECT 453.000 0.000 456.540 1.120 ;
  LAYER metal2 ;
  RECT 453.000 0.000 456.540 1.120 ;
  LAYER metal1 ;
  RECT 453.000 0.000 456.540 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 444.320 0.000 447.860 1.120 ;
  LAYER metal3 ;
  RECT 444.320 0.000 447.860 1.120 ;
  LAYER metal2 ;
  RECT 444.320 0.000 447.860 1.120 ;
  LAYER metal1 ;
  RECT 444.320 0.000 447.860 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER metal3 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER metal2 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER metal1 ;
  RECT 435.640 0.000 439.180 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 426.960 0.000 430.500 1.120 ;
  LAYER metal3 ;
  RECT 426.960 0.000 430.500 1.120 ;
  LAYER metal2 ;
  RECT 426.960 0.000 430.500 1.120 ;
  LAYER metal1 ;
  RECT 426.960 0.000 430.500 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 383.560 0.000 387.100 1.120 ;
  LAYER metal3 ;
  RECT 383.560 0.000 387.100 1.120 ;
  LAYER metal2 ;
  RECT 383.560 0.000 387.100 1.120 ;
  LAYER metal1 ;
  RECT 383.560 0.000 387.100 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 374.880 0.000 378.420 1.120 ;
  LAYER metal3 ;
  RECT 374.880 0.000 378.420 1.120 ;
  LAYER metal2 ;
  RECT 374.880 0.000 378.420 1.120 ;
  LAYER metal1 ;
  RECT 374.880 0.000 378.420 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 353.180 0.000 356.720 1.120 ;
  LAYER metal3 ;
  RECT 353.180 0.000 356.720 1.120 ;
  LAYER metal2 ;
  RECT 353.180 0.000 356.720 1.120 ;
  LAYER metal1 ;
  RECT 353.180 0.000 356.720 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER metal3 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER metal2 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER metal1 ;
  RECT 339.540 0.000 343.080 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 330.860 0.000 334.400 1.120 ;
  LAYER metal3 ;
  RECT 330.860 0.000 334.400 1.120 ;
  LAYER metal2 ;
  RECT 330.860 0.000 334.400 1.120 ;
  LAYER metal1 ;
  RECT 330.860 0.000 334.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 322.180 0.000 325.720 1.120 ;
  LAYER metal3 ;
  RECT 322.180 0.000 325.720 1.120 ;
  LAYER metal2 ;
  RECT 322.180 0.000 325.720 1.120 ;
  LAYER metal1 ;
  RECT 322.180 0.000 325.720 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 278.780 0.000 282.320 1.120 ;
  LAYER metal3 ;
  RECT 278.780 0.000 282.320 1.120 ;
  LAYER metal2 ;
  RECT 278.780 0.000 282.320 1.120 ;
  LAYER metal1 ;
  RECT 278.780 0.000 282.320 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 270.100 0.000 273.640 1.120 ;
  LAYER metal3 ;
  RECT 270.100 0.000 273.640 1.120 ;
  LAYER metal2 ;
  RECT 270.100 0.000 273.640 1.120 ;
  LAYER metal1 ;
  RECT 270.100 0.000 273.640 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER metal3 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER metal2 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER metal1 ;
  RECT 261.420 0.000 264.960 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER metal3 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER metal2 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER metal1 ;
  RECT 239.720 0.000 243.260 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 226.700 0.000 230.240 1.120 ;
  LAYER metal3 ;
  RECT 226.700 0.000 230.240 1.120 ;
  LAYER metal2 ;
  RECT 226.700 0.000 230.240 1.120 ;
  LAYER metal1 ;
  RECT 226.700 0.000 230.240 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 218.020 0.000 221.560 1.120 ;
  LAYER metal3 ;
  RECT 218.020 0.000 221.560 1.120 ;
  LAYER metal2 ;
  RECT 218.020 0.000 221.560 1.120 ;
  LAYER metal1 ;
  RECT 218.020 0.000 221.560 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 174.620 0.000 178.160 1.120 ;
  LAYER metal3 ;
  RECT 174.620 0.000 178.160 1.120 ;
  LAYER metal2 ;
  RECT 174.620 0.000 178.160 1.120 ;
  LAYER metal1 ;
  RECT 174.620 0.000 178.160 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 165.940 0.000 169.480 1.120 ;
  LAYER metal3 ;
  RECT 165.940 0.000 169.480 1.120 ;
  LAYER metal2 ;
  RECT 165.940 0.000 169.480 1.120 ;
  LAYER metal1 ;
  RECT 165.940 0.000 169.480 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 157.260 0.000 160.800 1.120 ;
  LAYER metal3 ;
  RECT 157.260 0.000 160.800 1.120 ;
  LAYER metal2 ;
  RECT 157.260 0.000 160.800 1.120 ;
  LAYER metal1 ;
  RECT 157.260 0.000 160.800 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 148.580 0.000 152.120 1.120 ;
  LAYER metal3 ;
  RECT 148.580 0.000 152.120 1.120 ;
  LAYER metal2 ;
  RECT 148.580 0.000 152.120 1.120 ;
  LAYER metal1 ;
  RECT 148.580 0.000 152.120 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER metal3 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER metal2 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER metal1 ;
  RECT 126.880 0.000 130.420 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal3 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal2 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal1 ;
  RECT 113.860 0.000 117.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal3 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal2 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal1 ;
  RECT 70.460 0.000 74.000 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 61.780 0.000 65.320 1.120 ;
  LAYER metal3 ;
  RECT 61.780 0.000 65.320 1.120 ;
  LAYER metal2 ;
  RECT 61.780 0.000 65.320 1.120 ;
  LAYER metal1 ;
  RECT 61.780 0.000 65.320 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 53.100 0.000 56.640 1.120 ;
  LAYER metal3 ;
  RECT 53.100 0.000 56.640 1.120 ;
  LAYER metal2 ;
  RECT 53.100 0.000 56.640 1.120 ;
  LAYER metal1 ;
  RECT 53.100 0.000 56.640 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 44.420 0.000 47.960 1.120 ;
  LAYER metal3 ;
  RECT 44.420 0.000 47.960 1.120 ;
  LAYER metal2 ;
  RECT 44.420 0.000 47.960 1.120 ;
  LAYER metal1 ;
  RECT 44.420 0.000 47.960 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal3 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal2 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal1 ;
  RECT 35.740 0.000 39.280 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal3 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal2 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal1 ;
  RECT 14.040 0.000 17.580 1.120 ;
 END
END VCC
PIN DO31
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1798.680 0.000 1799.800 1.120 ;
  LAYER metal3 ;
  RECT 1798.680 0.000 1799.800 1.120 ;
  LAYER metal2 ;
  RECT 1798.680 0.000 1799.800 1.120 ;
  LAYER metal1 ;
  RECT 1798.680 0.000 1799.800 1.120 ;
 END
END DO31
PIN DI31
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1790.620 0.000 1791.740 1.120 ;
  LAYER metal3 ;
  RECT 1790.620 0.000 1791.740 1.120 ;
  LAYER metal2 ;
  RECT 1790.620 0.000 1791.740 1.120 ;
  LAYER metal1 ;
  RECT 1790.620 0.000 1791.740 1.120 ;
 END
END DI31
PIN DO30
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1785.660 0.000 1786.780 1.120 ;
  LAYER metal3 ;
  RECT 1785.660 0.000 1786.780 1.120 ;
  LAYER metal2 ;
  RECT 1785.660 0.000 1786.780 1.120 ;
  LAYER metal1 ;
  RECT 1785.660 0.000 1786.780 1.120 ;
 END
END DO30
PIN DI30
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1776.980 0.000 1778.100 1.120 ;
  LAYER metal3 ;
  RECT 1776.980 0.000 1778.100 1.120 ;
  LAYER metal2 ;
  RECT 1776.980 0.000 1778.100 1.120 ;
  LAYER metal1 ;
  RECT 1776.980 0.000 1778.100 1.120 ;
 END
END DI30
PIN DO29
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1685.840 0.000 1686.960 1.120 ;
  LAYER metal3 ;
  RECT 1685.840 0.000 1686.960 1.120 ;
  LAYER metal2 ;
  RECT 1685.840 0.000 1686.960 1.120 ;
  LAYER metal1 ;
  RECT 1685.840 0.000 1686.960 1.120 ;
 END
END DO29
PIN DI29
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1677.160 0.000 1678.280 1.120 ;
  LAYER metal3 ;
  RECT 1677.160 0.000 1678.280 1.120 ;
  LAYER metal2 ;
  RECT 1677.160 0.000 1678.280 1.120 ;
  LAYER metal1 ;
  RECT 1677.160 0.000 1678.280 1.120 ;
 END
END DI29
PIN DO28
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1672.200 0.000 1673.320 1.120 ;
  LAYER metal3 ;
  RECT 1672.200 0.000 1673.320 1.120 ;
  LAYER metal2 ;
  RECT 1672.200 0.000 1673.320 1.120 ;
  LAYER metal1 ;
  RECT 1672.200 0.000 1673.320 1.120 ;
 END
END DO28
PIN DI28
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1664.140 0.000 1665.260 1.120 ;
  LAYER metal3 ;
  RECT 1664.140 0.000 1665.260 1.120 ;
  LAYER metal2 ;
  RECT 1664.140 0.000 1665.260 1.120 ;
  LAYER metal1 ;
  RECT 1664.140 0.000 1665.260 1.120 ;
 END
END DI28
PIN DO27
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1573.000 0.000 1574.120 1.120 ;
  LAYER metal3 ;
  RECT 1573.000 0.000 1574.120 1.120 ;
  LAYER metal2 ;
  RECT 1573.000 0.000 1574.120 1.120 ;
  LAYER metal1 ;
  RECT 1573.000 0.000 1574.120 1.120 ;
 END
END DO27
PIN DI27
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1564.320 0.000 1565.440 1.120 ;
  LAYER metal3 ;
  RECT 1564.320 0.000 1565.440 1.120 ;
  LAYER metal2 ;
  RECT 1564.320 0.000 1565.440 1.120 ;
  LAYER metal1 ;
  RECT 1564.320 0.000 1565.440 1.120 ;
 END
END DI27
PIN DO26
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1559.360 0.000 1560.480 1.120 ;
  LAYER metal3 ;
  RECT 1559.360 0.000 1560.480 1.120 ;
  LAYER metal2 ;
  RECT 1559.360 0.000 1560.480 1.120 ;
  LAYER metal1 ;
  RECT 1559.360 0.000 1560.480 1.120 ;
 END
END DO26
PIN DI26
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1551.300 0.000 1552.420 1.120 ;
  LAYER metal3 ;
  RECT 1551.300 0.000 1552.420 1.120 ;
  LAYER metal2 ;
  RECT 1551.300 0.000 1552.420 1.120 ;
  LAYER metal1 ;
  RECT 1551.300 0.000 1552.420 1.120 ;
 END
END DI26
PIN DO25
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1459.540 0.000 1460.660 1.120 ;
  LAYER metal3 ;
  RECT 1459.540 0.000 1460.660 1.120 ;
  LAYER metal2 ;
  RECT 1459.540 0.000 1460.660 1.120 ;
  LAYER metal1 ;
  RECT 1459.540 0.000 1460.660 1.120 ;
 END
END DO25
PIN DI25
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1451.480 0.000 1452.600 1.120 ;
  LAYER metal3 ;
  RECT 1451.480 0.000 1452.600 1.120 ;
  LAYER metal2 ;
  RECT 1451.480 0.000 1452.600 1.120 ;
  LAYER metal1 ;
  RECT 1451.480 0.000 1452.600 1.120 ;
 END
END DI25
PIN DO24
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1446.520 0.000 1447.640 1.120 ;
  LAYER metal3 ;
  RECT 1446.520 0.000 1447.640 1.120 ;
  LAYER metal2 ;
  RECT 1446.520 0.000 1447.640 1.120 ;
  LAYER metal1 ;
  RECT 1446.520 0.000 1447.640 1.120 ;
 END
END DO24
PIN DI24
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1437.840 0.000 1438.960 1.120 ;
  LAYER metal3 ;
  RECT 1437.840 0.000 1438.960 1.120 ;
  LAYER metal2 ;
  RECT 1437.840 0.000 1438.960 1.120 ;
  LAYER metal1 ;
  RECT 1437.840 0.000 1438.960 1.120 ;
 END
END DI24
PIN DO23
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1346.700 0.000 1347.820 1.120 ;
  LAYER metal3 ;
  RECT 1346.700 0.000 1347.820 1.120 ;
  LAYER metal2 ;
  RECT 1346.700 0.000 1347.820 1.120 ;
  LAYER metal1 ;
  RECT 1346.700 0.000 1347.820 1.120 ;
 END
END DO23
PIN DI23
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1338.020 0.000 1339.140 1.120 ;
  LAYER metal3 ;
  RECT 1338.020 0.000 1339.140 1.120 ;
  LAYER metal2 ;
  RECT 1338.020 0.000 1339.140 1.120 ;
  LAYER metal1 ;
  RECT 1338.020 0.000 1339.140 1.120 ;
 END
END DI23
PIN DO22
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1333.060 0.000 1334.180 1.120 ;
  LAYER metal3 ;
  RECT 1333.060 0.000 1334.180 1.120 ;
  LAYER metal2 ;
  RECT 1333.060 0.000 1334.180 1.120 ;
  LAYER metal1 ;
  RECT 1333.060 0.000 1334.180 1.120 ;
 END
END DO22
PIN DI22
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1325.000 0.000 1326.120 1.120 ;
  LAYER metal3 ;
  RECT 1325.000 0.000 1326.120 1.120 ;
  LAYER metal2 ;
  RECT 1325.000 0.000 1326.120 1.120 ;
  LAYER metal1 ;
  RECT 1325.000 0.000 1326.120 1.120 ;
 END
END DI22
PIN DO21
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1233.860 0.000 1234.980 1.120 ;
  LAYER metal3 ;
  RECT 1233.860 0.000 1234.980 1.120 ;
  LAYER metal2 ;
  RECT 1233.860 0.000 1234.980 1.120 ;
  LAYER metal1 ;
  RECT 1233.860 0.000 1234.980 1.120 ;
 END
END DO21
PIN DI21
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1225.180 0.000 1226.300 1.120 ;
  LAYER metal3 ;
  RECT 1225.180 0.000 1226.300 1.120 ;
  LAYER metal2 ;
  RECT 1225.180 0.000 1226.300 1.120 ;
  LAYER metal1 ;
  RECT 1225.180 0.000 1226.300 1.120 ;
 END
END DI21
PIN DO20
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1220.220 0.000 1221.340 1.120 ;
  LAYER metal3 ;
  RECT 1220.220 0.000 1221.340 1.120 ;
  LAYER metal2 ;
  RECT 1220.220 0.000 1221.340 1.120 ;
  LAYER metal1 ;
  RECT 1220.220 0.000 1221.340 1.120 ;
 END
END DO20
PIN DI20
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1212.160 0.000 1213.280 1.120 ;
  LAYER metal3 ;
  RECT 1212.160 0.000 1213.280 1.120 ;
  LAYER metal2 ;
  RECT 1212.160 0.000 1213.280 1.120 ;
  LAYER metal1 ;
  RECT 1212.160 0.000 1213.280 1.120 ;
 END
END DI20
PIN DO19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1120.400 0.000 1121.520 1.120 ;
  LAYER metal3 ;
  RECT 1120.400 0.000 1121.520 1.120 ;
  LAYER metal2 ;
  RECT 1120.400 0.000 1121.520 1.120 ;
  LAYER metal1 ;
  RECT 1120.400 0.000 1121.520 1.120 ;
 END
END DO19
PIN DI19
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1112.340 0.000 1113.460 1.120 ;
  LAYER metal3 ;
  RECT 1112.340 0.000 1113.460 1.120 ;
  LAYER metal2 ;
  RECT 1112.340 0.000 1113.460 1.120 ;
  LAYER metal1 ;
  RECT 1112.340 0.000 1113.460 1.120 ;
 END
END DI19
PIN DO18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1107.380 0.000 1108.500 1.120 ;
  LAYER metal3 ;
  RECT 1107.380 0.000 1108.500 1.120 ;
  LAYER metal2 ;
  RECT 1107.380 0.000 1108.500 1.120 ;
  LAYER metal1 ;
  RECT 1107.380 0.000 1108.500 1.120 ;
 END
END DO18
PIN DI18
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 1098.700 0.000 1099.820 1.120 ;
  LAYER metal3 ;
  RECT 1098.700 0.000 1099.820 1.120 ;
  LAYER metal2 ;
  RECT 1098.700 0.000 1099.820 1.120 ;
  LAYER metal1 ;
  RECT 1098.700 0.000 1099.820 1.120 ;
 END
END DI18
PIN DO17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 1007.560 0.000 1008.680 1.120 ;
  LAYER metal3 ;
  RECT 1007.560 0.000 1008.680 1.120 ;
  LAYER metal2 ;
  RECT 1007.560 0.000 1008.680 1.120 ;
  LAYER metal1 ;
  RECT 1007.560 0.000 1008.680 1.120 ;
 END
END DO17
PIN DI17
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 998.880 0.000 1000.000 1.120 ;
  LAYER metal3 ;
  RECT 998.880 0.000 1000.000 1.120 ;
  LAYER metal2 ;
  RECT 998.880 0.000 1000.000 1.120 ;
  LAYER metal1 ;
  RECT 998.880 0.000 1000.000 1.120 ;
 END
END DI17
PIN DO16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 994.540 0.000 995.660 1.120 ;
  LAYER metal3 ;
  RECT 994.540 0.000 995.660 1.120 ;
  LAYER metal2 ;
  RECT 994.540 0.000 995.660 1.120 ;
  LAYER metal1 ;
  RECT 994.540 0.000 995.660 1.120 ;
 END
END DO16
PIN DI16
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 985.860 0.000 986.980 1.120 ;
  LAYER metal3 ;
  RECT 985.860 0.000 986.980 1.120 ;
  LAYER metal2 ;
  RECT 985.860 0.000 986.980 1.120 ;
  LAYER metal1 ;
  RECT 985.860 0.000 986.980 1.120 ;
 END
END DI16
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 980.280 0.000 981.400 1.120 ;
  LAYER metal3 ;
  RECT 980.280 0.000 981.400 1.120 ;
  LAYER metal2 ;
  RECT 980.280 0.000 981.400 1.120 ;
  LAYER metal1 ;
  RECT 980.280 0.000 981.400 1.120 ;
 END
END A1
PIN WEB
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 978.420 0.000 979.540 1.120 ;
  LAYER metal3 ;
  RECT 978.420 0.000 979.540 1.120 ;
  LAYER metal2 ;
  RECT 978.420 0.000 979.540 1.120 ;
  LAYER metal1 ;
  RECT 978.420 0.000 979.540 1.120 ;
 END
END WEB
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.033 ;
 PORT
  LAYER metal4 ;
  RECT 973.460 0.000 974.580 1.120 ;
  LAYER metal3 ;
  RECT 973.460 0.000 974.580 1.120 ;
  LAYER metal2 ;
  RECT 973.460 0.000 974.580 1.120 ;
  LAYER metal1 ;
  RECT 973.460 0.000 974.580 1.120 ;
 END
END OE
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.123 ;
 PORT
  LAYER metal4 ;
  RECT 971.600 0.000 972.720 1.120 ;
  LAYER metal3 ;
  RECT 971.600 0.000 972.720 1.120 ;
  LAYER metal2 ;
  RECT 971.600 0.000 972.720 1.120 ;
  LAYER metal1 ;
  RECT 971.600 0.000 972.720 1.120 ;
 END
END CS
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 969.740 0.000 970.860 1.120 ;
  LAYER metal3 ;
  RECT 969.740 0.000 970.860 1.120 ;
  LAYER metal2 ;
  RECT 969.740 0.000 970.860 1.120 ;
  LAYER metal1 ;
  RECT 969.740 0.000 970.860 1.120 ;
 END
END A3
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 962.920 0.000 964.040 1.120 ;
  LAYER metal3 ;
  RECT 962.920 0.000 964.040 1.120 ;
  LAYER metal2 ;
  RECT 962.920 0.000 964.040 1.120 ;
  LAYER metal1 ;
  RECT 962.920 0.000 964.040 1.120 ;
 END
END A4
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 949.900 0.000 951.020 1.120 ;
  LAYER metal3 ;
  RECT 949.900 0.000 951.020 1.120 ;
  LAYER metal2 ;
  RECT 949.900 0.000 951.020 1.120 ;
  LAYER metal1 ;
  RECT 949.900 0.000 951.020 1.120 ;
 END
END A2
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.063 ;
 PORT
  LAYER metal4 ;
  RECT 946.800 0.000 947.920 1.120 ;
  LAYER metal3 ;
  RECT 946.800 0.000 947.920 1.120 ;
  LAYER metal2 ;
  RECT 946.800 0.000 947.920 1.120 ;
  LAYER metal1 ;
  RECT 946.800 0.000 947.920 1.120 ;
 END
END CK
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 944.940 0.000 946.060 1.120 ;
  LAYER metal3 ;
  RECT 944.940 0.000 946.060 1.120 ;
  LAYER metal2 ;
  RECT 944.940 0.000 946.060 1.120 ;
  LAYER metal1 ;
  RECT 944.940 0.000 946.060 1.120 ;
 END
END A0
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 940.600 0.000 941.720 1.120 ;
  LAYER metal3 ;
  RECT 940.600 0.000 941.720 1.120 ;
  LAYER metal2 ;
  RECT 940.600 0.000 941.720 1.120 ;
  LAYER metal1 ;
  RECT 940.600 0.000 941.720 1.120 ;
 END
END A5
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 933.160 0.000 934.280 1.120 ;
  LAYER metal3 ;
  RECT 933.160 0.000 934.280 1.120 ;
  LAYER metal2 ;
  RECT 933.160 0.000 934.280 1.120 ;
  LAYER metal1 ;
  RECT 933.160 0.000 934.280 1.120 ;
 END
END A6
PIN A7
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 930.060 0.000 931.180 1.120 ;
  LAYER metal3 ;
  RECT 930.060 0.000 931.180 1.120 ;
  LAYER metal2 ;
  RECT 930.060 0.000 931.180 1.120 ;
  LAYER metal1 ;
  RECT 930.060 0.000 931.180 1.120 ;
 END
END A7
PIN A8
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 922.000 0.000 923.120 1.120 ;
  LAYER metal3 ;
  RECT 922.000 0.000 923.120 1.120 ;
  LAYER metal2 ;
  RECT 922.000 0.000 923.120 1.120 ;
  LAYER metal1 ;
  RECT 922.000 0.000 923.120 1.120 ;
 END
END A8
PIN DO15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 824.660 0.000 825.780 1.120 ;
  LAYER metal3 ;
  RECT 824.660 0.000 825.780 1.120 ;
  LAYER metal2 ;
  RECT 824.660 0.000 825.780 1.120 ;
  LAYER metal1 ;
  RECT 824.660 0.000 825.780 1.120 ;
 END
END DO15
PIN DI15
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 815.980 0.000 817.100 1.120 ;
  LAYER metal3 ;
  RECT 815.980 0.000 817.100 1.120 ;
  LAYER metal2 ;
  RECT 815.980 0.000 817.100 1.120 ;
  LAYER metal1 ;
  RECT 815.980 0.000 817.100 1.120 ;
 END
END DI15
PIN DO14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 811.640 0.000 812.760 1.120 ;
  LAYER metal3 ;
  RECT 811.640 0.000 812.760 1.120 ;
  LAYER metal2 ;
  RECT 811.640 0.000 812.760 1.120 ;
  LAYER metal1 ;
  RECT 811.640 0.000 812.760 1.120 ;
 END
END DO14
PIN DI14
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 802.960 0.000 804.080 1.120 ;
  LAYER metal3 ;
  RECT 802.960 0.000 804.080 1.120 ;
  LAYER metal2 ;
  RECT 802.960 0.000 804.080 1.120 ;
  LAYER metal1 ;
  RECT 802.960 0.000 804.080 1.120 ;
 END
END DI14
PIN DO13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 711.820 0.000 712.940 1.120 ;
  LAYER metal3 ;
  RECT 711.820 0.000 712.940 1.120 ;
  LAYER metal2 ;
  RECT 711.820 0.000 712.940 1.120 ;
  LAYER metal1 ;
  RECT 711.820 0.000 712.940 1.120 ;
 END
END DO13
PIN DI13
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 703.140 0.000 704.260 1.120 ;
  LAYER metal3 ;
  RECT 703.140 0.000 704.260 1.120 ;
  LAYER metal2 ;
  RECT 703.140 0.000 704.260 1.120 ;
  LAYER metal1 ;
  RECT 703.140 0.000 704.260 1.120 ;
 END
END DI13
PIN DO12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 698.180 0.000 699.300 1.120 ;
  LAYER metal3 ;
  RECT 698.180 0.000 699.300 1.120 ;
  LAYER metal2 ;
  RECT 698.180 0.000 699.300 1.120 ;
  LAYER metal1 ;
  RECT 698.180 0.000 699.300 1.120 ;
 END
END DO12
PIN DI12
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 690.120 0.000 691.240 1.120 ;
  LAYER metal3 ;
  RECT 690.120 0.000 691.240 1.120 ;
  LAYER metal2 ;
  RECT 690.120 0.000 691.240 1.120 ;
  LAYER metal1 ;
  RECT 690.120 0.000 691.240 1.120 ;
 END
END DI12
PIN DO11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 598.360 0.000 599.480 1.120 ;
  LAYER metal3 ;
  RECT 598.360 0.000 599.480 1.120 ;
  LAYER metal2 ;
  RECT 598.360 0.000 599.480 1.120 ;
  LAYER metal1 ;
  RECT 598.360 0.000 599.480 1.120 ;
 END
END DO11
PIN DI11
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 590.300 0.000 591.420 1.120 ;
  LAYER metal3 ;
  RECT 590.300 0.000 591.420 1.120 ;
  LAYER metal2 ;
  RECT 590.300 0.000 591.420 1.120 ;
  LAYER metal1 ;
  RECT 590.300 0.000 591.420 1.120 ;
 END
END DI11
PIN DO10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 585.340 0.000 586.460 1.120 ;
  LAYER metal3 ;
  RECT 585.340 0.000 586.460 1.120 ;
  LAYER metal2 ;
  RECT 585.340 0.000 586.460 1.120 ;
  LAYER metal1 ;
  RECT 585.340 0.000 586.460 1.120 ;
 END
END DO10
PIN DI10
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 576.660 0.000 577.780 1.120 ;
  LAYER metal3 ;
  RECT 576.660 0.000 577.780 1.120 ;
  LAYER metal2 ;
  RECT 576.660 0.000 577.780 1.120 ;
  LAYER metal1 ;
  RECT 576.660 0.000 577.780 1.120 ;
 END
END DI10
PIN DO9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 485.520 0.000 486.640 1.120 ;
  LAYER metal3 ;
  RECT 485.520 0.000 486.640 1.120 ;
  LAYER metal2 ;
  RECT 485.520 0.000 486.640 1.120 ;
  LAYER metal1 ;
  RECT 485.520 0.000 486.640 1.120 ;
 END
END DO9
PIN DI9
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 476.840 0.000 477.960 1.120 ;
  LAYER metal3 ;
  RECT 476.840 0.000 477.960 1.120 ;
  LAYER metal2 ;
  RECT 476.840 0.000 477.960 1.120 ;
  LAYER metal1 ;
  RECT 476.840 0.000 477.960 1.120 ;
 END
END DI9
PIN DO8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 472.500 0.000 473.620 1.120 ;
  LAYER metal3 ;
  RECT 472.500 0.000 473.620 1.120 ;
  LAYER metal2 ;
  RECT 472.500 0.000 473.620 1.120 ;
  LAYER metal1 ;
  RECT 472.500 0.000 473.620 1.120 ;
 END
END DO8
PIN DI8
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 463.820 0.000 464.940 1.120 ;
  LAYER metal3 ;
  RECT 463.820 0.000 464.940 1.120 ;
  LAYER metal2 ;
  RECT 463.820 0.000 464.940 1.120 ;
  LAYER metal1 ;
  RECT 463.820 0.000 464.940 1.120 ;
 END
END DI8
PIN DO7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 372.680 0.000 373.800 1.120 ;
  LAYER metal3 ;
  RECT 372.680 0.000 373.800 1.120 ;
  LAYER metal2 ;
  RECT 372.680 0.000 373.800 1.120 ;
  LAYER metal1 ;
  RECT 372.680 0.000 373.800 1.120 ;
 END
END DO7
PIN DI7
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 364.000 0.000 365.120 1.120 ;
  LAYER metal3 ;
  RECT 364.000 0.000 365.120 1.120 ;
  LAYER metal2 ;
  RECT 364.000 0.000 365.120 1.120 ;
  LAYER metal1 ;
  RECT 364.000 0.000 365.120 1.120 ;
 END
END DI7
PIN DO6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER metal3 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER metal2 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER metal1 ;
  RECT 359.040 0.000 360.160 1.120 ;
 END
END DO6
PIN DI6
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 350.980 0.000 352.100 1.120 ;
  LAYER metal3 ;
  RECT 350.980 0.000 352.100 1.120 ;
  LAYER metal2 ;
  RECT 350.980 0.000 352.100 1.120 ;
  LAYER metal1 ;
  RECT 350.980 0.000 352.100 1.120 ;
 END
END DI6
PIN DO5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER metal3 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER metal2 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER metal1 ;
  RECT 259.220 0.000 260.340 1.120 ;
 END
END DO5
PIN DI5
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER metal3 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER metal2 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER metal1 ;
  RECT 251.160 0.000 252.280 1.120 ;
 END
END DI5
PIN DO4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER metal3 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER metal2 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER metal1 ;
  RECT 246.200 0.000 247.320 1.120 ;
 END
END DO4
PIN DI4
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER metal3 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER metal2 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER metal1 ;
  RECT 237.520 0.000 238.640 1.120 ;
 END
END DI4
PIN DO3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal3 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal2 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal1 ;
  RECT 146.380 0.000 147.500 1.120 ;
 END
END DO3
PIN DI3
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER metal3 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER metal2 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER metal1 ;
  RECT 137.700 0.000 138.820 1.120 ;
 END
END DI3
PIN DO2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER metal3 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER metal2 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER metal1 ;
  RECT 133.360 0.000 134.480 1.120 ;
 END
END DO2
PIN DI2
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER metal3 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER metal2 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER metal1 ;
  RECT 124.680 0.000 125.800 1.120 ;
 END
END DI2
PIN DO1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal3 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal2 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal1 ;
  RECT 33.540 0.000 34.660 1.120 ;
 END
END DO1
PIN DI1
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal3 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal2 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal1 ;
  RECT 24.860 0.000 25.980 1.120 ;
 END
END DI1
PIN DO0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.116 ;
 PORT
  LAYER metal4 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal3 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal2 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal1 ;
  RECT 19.900 0.000 21.020 1.120 ;
 END
END DO0
PIN DI0
  DIRECTION INPUT ;
  CAPACITANCE 0.039 ;
 PORT
  LAYER metal4 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal3 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal2 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal1 ;
  RECT 11.840 0.000 12.960 1.120 ;
 END
END DI0
OBS
  LAYER metal1 SPACING 0.280 ;
  RECT 0.000 0.140 1899.060 166.880 ;
  LAYER metal2 SPACING 0.320 ;
  RECT 0.000 0.140 1899.060 166.880 ;
  LAYER metal3 SPACING 0.320 ;
  RECT 0.000 0.140 1899.060 166.880 ;
  LAYER metal4 SPACING 0.600 ;
  RECT 0.000 0.140 1899.060 166.880 ;
  LAYER via ;
  RECT 0.000 0.140 1899.060 166.880 ;
  LAYER via2 ;
  RECT 0.000 0.140 1899.060 166.880 ;
  LAYER via3 ;
  RECT 0.000 0.140 1899.060 166.880 ;
END
END SUMA180_384X32X1BM4
END LIBRARY



