# 
#              Synchronous Dual Port SRAM Compiler 
# 
#                    UMC 0.18um Generic Logic Process 
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : SJMA180_32768X16X1BM8
#       Words            : 32768
#       Bits             : 16
#       Byte-Write       : 1
#       Aspect Ratio     : 8
#       Output Loading   : 0.5  (pf)
#       Data Slew        : 0.5  (ns)
#       CK Slew          : 0.5  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2022/01/19 09:49:47
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO SJMA180_32768X16X1BM8
CLASS BLOCK ;
FOREIGN SJMA180_32768X16X1BM8 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 3613.980 BY 1711.920 ;
SYMMETRY x y r90 ;
SITE core ;
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal5 ;
  RECT 3612.860 1697.140 3613.980 1700.380 ;
  LAYER metal4 ;
  RECT 3612.860 1697.140 3613.980 1700.380 ;
  LAYER metal3 ;
  RECT 3612.860 1697.140 3613.980 1700.380 ;
  LAYER metal2 ;
  RECT 3612.860 1697.140 3613.980 1700.380 ;
  LAYER metal1 ;
  RECT 3612.860 1697.140 3613.980 1700.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1689.300 3613.980 1692.540 ;
  LAYER metal4 ;
  RECT 3612.860 1689.300 3613.980 1692.540 ;
  LAYER metal3 ;
  RECT 3612.860 1689.300 3613.980 1692.540 ;
  LAYER metal2 ;
  RECT 3612.860 1689.300 3613.980 1692.540 ;
  LAYER metal1 ;
  RECT 3612.860 1689.300 3613.980 1692.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1681.460 3613.980 1684.700 ;
  LAYER metal4 ;
  RECT 3612.860 1681.460 3613.980 1684.700 ;
  LAYER metal3 ;
  RECT 3612.860 1681.460 3613.980 1684.700 ;
  LAYER metal2 ;
  RECT 3612.860 1681.460 3613.980 1684.700 ;
  LAYER metal1 ;
  RECT 3612.860 1681.460 3613.980 1684.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1673.620 3613.980 1676.860 ;
  LAYER metal4 ;
  RECT 3612.860 1673.620 3613.980 1676.860 ;
  LAYER metal3 ;
  RECT 3612.860 1673.620 3613.980 1676.860 ;
  LAYER metal2 ;
  RECT 3612.860 1673.620 3613.980 1676.860 ;
  LAYER metal1 ;
  RECT 3612.860 1673.620 3613.980 1676.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1665.780 3613.980 1669.020 ;
  LAYER metal4 ;
  RECT 3612.860 1665.780 3613.980 1669.020 ;
  LAYER metal3 ;
  RECT 3612.860 1665.780 3613.980 1669.020 ;
  LAYER metal2 ;
  RECT 3612.860 1665.780 3613.980 1669.020 ;
  LAYER metal1 ;
  RECT 3612.860 1665.780 3613.980 1669.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1657.940 3613.980 1661.180 ;
  LAYER metal4 ;
  RECT 3612.860 1657.940 3613.980 1661.180 ;
  LAYER metal3 ;
  RECT 3612.860 1657.940 3613.980 1661.180 ;
  LAYER metal2 ;
  RECT 3612.860 1657.940 3613.980 1661.180 ;
  LAYER metal1 ;
  RECT 3612.860 1657.940 3613.980 1661.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1618.740 3613.980 1621.980 ;
  LAYER metal4 ;
  RECT 3612.860 1618.740 3613.980 1621.980 ;
  LAYER metal3 ;
  RECT 3612.860 1618.740 3613.980 1621.980 ;
  LAYER metal2 ;
  RECT 3612.860 1618.740 3613.980 1621.980 ;
  LAYER metal1 ;
  RECT 3612.860 1618.740 3613.980 1621.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1610.900 3613.980 1614.140 ;
  LAYER metal4 ;
  RECT 3612.860 1610.900 3613.980 1614.140 ;
  LAYER metal3 ;
  RECT 3612.860 1610.900 3613.980 1614.140 ;
  LAYER metal2 ;
  RECT 3612.860 1610.900 3613.980 1614.140 ;
  LAYER metal1 ;
  RECT 3612.860 1610.900 3613.980 1614.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1603.060 3613.980 1606.300 ;
  LAYER metal4 ;
  RECT 3612.860 1603.060 3613.980 1606.300 ;
  LAYER metal3 ;
  RECT 3612.860 1603.060 3613.980 1606.300 ;
  LAYER metal2 ;
  RECT 3612.860 1603.060 3613.980 1606.300 ;
  LAYER metal1 ;
  RECT 3612.860 1603.060 3613.980 1606.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1595.220 3613.980 1598.460 ;
  LAYER metal4 ;
  RECT 3612.860 1595.220 3613.980 1598.460 ;
  LAYER metal3 ;
  RECT 3612.860 1595.220 3613.980 1598.460 ;
  LAYER metal2 ;
  RECT 3612.860 1595.220 3613.980 1598.460 ;
  LAYER metal1 ;
  RECT 3612.860 1595.220 3613.980 1598.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1587.380 3613.980 1590.620 ;
  LAYER metal4 ;
  RECT 3612.860 1587.380 3613.980 1590.620 ;
  LAYER metal3 ;
  RECT 3612.860 1587.380 3613.980 1590.620 ;
  LAYER metal2 ;
  RECT 3612.860 1587.380 3613.980 1590.620 ;
  LAYER metal1 ;
  RECT 3612.860 1587.380 3613.980 1590.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1579.540 3613.980 1582.780 ;
  LAYER metal4 ;
  RECT 3612.860 1579.540 3613.980 1582.780 ;
  LAYER metal3 ;
  RECT 3612.860 1579.540 3613.980 1582.780 ;
  LAYER metal2 ;
  RECT 3612.860 1579.540 3613.980 1582.780 ;
  LAYER metal1 ;
  RECT 3612.860 1579.540 3613.980 1582.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1540.340 3613.980 1543.580 ;
  LAYER metal4 ;
  RECT 3612.860 1540.340 3613.980 1543.580 ;
  LAYER metal3 ;
  RECT 3612.860 1540.340 3613.980 1543.580 ;
  LAYER metal2 ;
  RECT 3612.860 1540.340 3613.980 1543.580 ;
  LAYER metal1 ;
  RECT 3612.860 1540.340 3613.980 1543.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1532.500 3613.980 1535.740 ;
  LAYER metal4 ;
  RECT 3612.860 1532.500 3613.980 1535.740 ;
  LAYER metal3 ;
  RECT 3612.860 1532.500 3613.980 1535.740 ;
  LAYER metal2 ;
  RECT 3612.860 1532.500 3613.980 1535.740 ;
  LAYER metal1 ;
  RECT 3612.860 1532.500 3613.980 1535.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1524.660 3613.980 1527.900 ;
  LAYER metal4 ;
  RECT 3612.860 1524.660 3613.980 1527.900 ;
  LAYER metal3 ;
  RECT 3612.860 1524.660 3613.980 1527.900 ;
  LAYER metal2 ;
  RECT 3612.860 1524.660 3613.980 1527.900 ;
  LAYER metal1 ;
  RECT 3612.860 1524.660 3613.980 1527.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1516.820 3613.980 1520.060 ;
  LAYER metal4 ;
  RECT 3612.860 1516.820 3613.980 1520.060 ;
  LAYER metal3 ;
  RECT 3612.860 1516.820 3613.980 1520.060 ;
  LAYER metal2 ;
  RECT 3612.860 1516.820 3613.980 1520.060 ;
  LAYER metal1 ;
  RECT 3612.860 1516.820 3613.980 1520.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1508.980 3613.980 1512.220 ;
  LAYER metal4 ;
  RECT 3612.860 1508.980 3613.980 1512.220 ;
  LAYER metal3 ;
  RECT 3612.860 1508.980 3613.980 1512.220 ;
  LAYER metal2 ;
  RECT 3612.860 1508.980 3613.980 1512.220 ;
  LAYER metal1 ;
  RECT 3612.860 1508.980 3613.980 1512.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1501.140 3613.980 1504.380 ;
  LAYER metal4 ;
  RECT 3612.860 1501.140 3613.980 1504.380 ;
  LAYER metal3 ;
  RECT 3612.860 1501.140 3613.980 1504.380 ;
  LAYER metal2 ;
  RECT 3612.860 1501.140 3613.980 1504.380 ;
  LAYER metal1 ;
  RECT 3612.860 1501.140 3613.980 1504.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1461.940 3613.980 1465.180 ;
  LAYER metal4 ;
  RECT 3612.860 1461.940 3613.980 1465.180 ;
  LAYER metal3 ;
  RECT 3612.860 1461.940 3613.980 1465.180 ;
  LAYER metal2 ;
  RECT 3612.860 1461.940 3613.980 1465.180 ;
  LAYER metal1 ;
  RECT 3612.860 1461.940 3613.980 1465.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1454.100 3613.980 1457.340 ;
  LAYER metal4 ;
  RECT 3612.860 1454.100 3613.980 1457.340 ;
  LAYER metal3 ;
  RECT 3612.860 1454.100 3613.980 1457.340 ;
  LAYER metal2 ;
  RECT 3612.860 1454.100 3613.980 1457.340 ;
  LAYER metal1 ;
  RECT 3612.860 1454.100 3613.980 1457.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1446.260 3613.980 1449.500 ;
  LAYER metal4 ;
  RECT 3612.860 1446.260 3613.980 1449.500 ;
  LAYER metal3 ;
  RECT 3612.860 1446.260 3613.980 1449.500 ;
  LAYER metal2 ;
  RECT 3612.860 1446.260 3613.980 1449.500 ;
  LAYER metal1 ;
  RECT 3612.860 1446.260 3613.980 1449.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1438.420 3613.980 1441.660 ;
  LAYER metal4 ;
  RECT 3612.860 1438.420 3613.980 1441.660 ;
  LAYER metal3 ;
  RECT 3612.860 1438.420 3613.980 1441.660 ;
  LAYER metal2 ;
  RECT 3612.860 1438.420 3613.980 1441.660 ;
  LAYER metal1 ;
  RECT 3612.860 1438.420 3613.980 1441.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1430.580 3613.980 1433.820 ;
  LAYER metal4 ;
  RECT 3612.860 1430.580 3613.980 1433.820 ;
  LAYER metal3 ;
  RECT 3612.860 1430.580 3613.980 1433.820 ;
  LAYER metal2 ;
  RECT 3612.860 1430.580 3613.980 1433.820 ;
  LAYER metal1 ;
  RECT 3612.860 1430.580 3613.980 1433.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1422.740 3613.980 1425.980 ;
  LAYER metal4 ;
  RECT 3612.860 1422.740 3613.980 1425.980 ;
  LAYER metal3 ;
  RECT 3612.860 1422.740 3613.980 1425.980 ;
  LAYER metal2 ;
  RECT 3612.860 1422.740 3613.980 1425.980 ;
  LAYER metal1 ;
  RECT 3612.860 1422.740 3613.980 1425.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1383.540 3613.980 1386.780 ;
  LAYER metal4 ;
  RECT 3612.860 1383.540 3613.980 1386.780 ;
  LAYER metal3 ;
  RECT 3612.860 1383.540 3613.980 1386.780 ;
  LAYER metal2 ;
  RECT 3612.860 1383.540 3613.980 1386.780 ;
  LAYER metal1 ;
  RECT 3612.860 1383.540 3613.980 1386.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1375.700 3613.980 1378.940 ;
  LAYER metal4 ;
  RECT 3612.860 1375.700 3613.980 1378.940 ;
  LAYER metal3 ;
  RECT 3612.860 1375.700 3613.980 1378.940 ;
  LAYER metal2 ;
  RECT 3612.860 1375.700 3613.980 1378.940 ;
  LAYER metal1 ;
  RECT 3612.860 1375.700 3613.980 1378.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1367.860 3613.980 1371.100 ;
  LAYER metal4 ;
  RECT 3612.860 1367.860 3613.980 1371.100 ;
  LAYER metal3 ;
  RECT 3612.860 1367.860 3613.980 1371.100 ;
  LAYER metal2 ;
  RECT 3612.860 1367.860 3613.980 1371.100 ;
  LAYER metal1 ;
  RECT 3612.860 1367.860 3613.980 1371.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1360.020 3613.980 1363.260 ;
  LAYER metal4 ;
  RECT 3612.860 1360.020 3613.980 1363.260 ;
  LAYER metal3 ;
  RECT 3612.860 1360.020 3613.980 1363.260 ;
  LAYER metal2 ;
  RECT 3612.860 1360.020 3613.980 1363.260 ;
  LAYER metal1 ;
  RECT 3612.860 1360.020 3613.980 1363.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1352.180 3613.980 1355.420 ;
  LAYER metal4 ;
  RECT 3612.860 1352.180 3613.980 1355.420 ;
  LAYER metal3 ;
  RECT 3612.860 1352.180 3613.980 1355.420 ;
  LAYER metal2 ;
  RECT 3612.860 1352.180 3613.980 1355.420 ;
  LAYER metal1 ;
  RECT 3612.860 1352.180 3613.980 1355.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1344.340 3613.980 1347.580 ;
  LAYER metal4 ;
  RECT 3612.860 1344.340 3613.980 1347.580 ;
  LAYER metal3 ;
  RECT 3612.860 1344.340 3613.980 1347.580 ;
  LAYER metal2 ;
  RECT 3612.860 1344.340 3613.980 1347.580 ;
  LAYER metal1 ;
  RECT 3612.860 1344.340 3613.980 1347.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1305.140 3613.980 1308.380 ;
  LAYER metal4 ;
  RECT 3612.860 1305.140 3613.980 1308.380 ;
  LAYER metal3 ;
  RECT 3612.860 1305.140 3613.980 1308.380 ;
  LAYER metal2 ;
  RECT 3612.860 1305.140 3613.980 1308.380 ;
  LAYER metal1 ;
  RECT 3612.860 1305.140 3613.980 1308.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1297.300 3613.980 1300.540 ;
  LAYER metal4 ;
  RECT 3612.860 1297.300 3613.980 1300.540 ;
  LAYER metal3 ;
  RECT 3612.860 1297.300 3613.980 1300.540 ;
  LAYER metal2 ;
  RECT 3612.860 1297.300 3613.980 1300.540 ;
  LAYER metal1 ;
  RECT 3612.860 1297.300 3613.980 1300.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1289.460 3613.980 1292.700 ;
  LAYER metal4 ;
  RECT 3612.860 1289.460 3613.980 1292.700 ;
  LAYER metal3 ;
  RECT 3612.860 1289.460 3613.980 1292.700 ;
  LAYER metal2 ;
  RECT 3612.860 1289.460 3613.980 1292.700 ;
  LAYER metal1 ;
  RECT 3612.860 1289.460 3613.980 1292.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1281.620 3613.980 1284.860 ;
  LAYER metal4 ;
  RECT 3612.860 1281.620 3613.980 1284.860 ;
  LAYER metal3 ;
  RECT 3612.860 1281.620 3613.980 1284.860 ;
  LAYER metal2 ;
  RECT 3612.860 1281.620 3613.980 1284.860 ;
  LAYER metal1 ;
  RECT 3612.860 1281.620 3613.980 1284.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1273.780 3613.980 1277.020 ;
  LAYER metal4 ;
  RECT 3612.860 1273.780 3613.980 1277.020 ;
  LAYER metal3 ;
  RECT 3612.860 1273.780 3613.980 1277.020 ;
  LAYER metal2 ;
  RECT 3612.860 1273.780 3613.980 1277.020 ;
  LAYER metal1 ;
  RECT 3612.860 1273.780 3613.980 1277.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1265.940 3613.980 1269.180 ;
  LAYER metal4 ;
  RECT 3612.860 1265.940 3613.980 1269.180 ;
  LAYER metal3 ;
  RECT 3612.860 1265.940 3613.980 1269.180 ;
  LAYER metal2 ;
  RECT 3612.860 1265.940 3613.980 1269.180 ;
  LAYER metal1 ;
  RECT 3612.860 1265.940 3613.980 1269.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1226.740 3613.980 1229.980 ;
  LAYER metal4 ;
  RECT 3612.860 1226.740 3613.980 1229.980 ;
  LAYER metal3 ;
  RECT 3612.860 1226.740 3613.980 1229.980 ;
  LAYER metal2 ;
  RECT 3612.860 1226.740 3613.980 1229.980 ;
  LAYER metal1 ;
  RECT 3612.860 1226.740 3613.980 1229.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1218.900 3613.980 1222.140 ;
  LAYER metal4 ;
  RECT 3612.860 1218.900 3613.980 1222.140 ;
  LAYER metal3 ;
  RECT 3612.860 1218.900 3613.980 1222.140 ;
  LAYER metal2 ;
  RECT 3612.860 1218.900 3613.980 1222.140 ;
  LAYER metal1 ;
  RECT 3612.860 1218.900 3613.980 1222.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1211.060 3613.980 1214.300 ;
  LAYER metal4 ;
  RECT 3612.860 1211.060 3613.980 1214.300 ;
  LAYER metal3 ;
  RECT 3612.860 1211.060 3613.980 1214.300 ;
  LAYER metal2 ;
  RECT 3612.860 1211.060 3613.980 1214.300 ;
  LAYER metal1 ;
  RECT 3612.860 1211.060 3613.980 1214.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1203.220 3613.980 1206.460 ;
  LAYER metal4 ;
  RECT 3612.860 1203.220 3613.980 1206.460 ;
  LAYER metal3 ;
  RECT 3612.860 1203.220 3613.980 1206.460 ;
  LAYER metal2 ;
  RECT 3612.860 1203.220 3613.980 1206.460 ;
  LAYER metal1 ;
  RECT 3612.860 1203.220 3613.980 1206.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1195.380 3613.980 1198.620 ;
  LAYER metal4 ;
  RECT 3612.860 1195.380 3613.980 1198.620 ;
  LAYER metal3 ;
  RECT 3612.860 1195.380 3613.980 1198.620 ;
  LAYER metal2 ;
  RECT 3612.860 1195.380 3613.980 1198.620 ;
  LAYER metal1 ;
  RECT 3612.860 1195.380 3613.980 1198.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1187.540 3613.980 1190.780 ;
  LAYER metal4 ;
  RECT 3612.860 1187.540 3613.980 1190.780 ;
  LAYER metal3 ;
  RECT 3612.860 1187.540 3613.980 1190.780 ;
  LAYER metal2 ;
  RECT 3612.860 1187.540 3613.980 1190.780 ;
  LAYER metal1 ;
  RECT 3612.860 1187.540 3613.980 1190.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1148.340 3613.980 1151.580 ;
  LAYER metal4 ;
  RECT 3612.860 1148.340 3613.980 1151.580 ;
  LAYER metal3 ;
  RECT 3612.860 1148.340 3613.980 1151.580 ;
  LAYER metal2 ;
  RECT 3612.860 1148.340 3613.980 1151.580 ;
  LAYER metal1 ;
  RECT 3612.860 1148.340 3613.980 1151.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1140.500 3613.980 1143.740 ;
  LAYER metal4 ;
  RECT 3612.860 1140.500 3613.980 1143.740 ;
  LAYER metal3 ;
  RECT 3612.860 1140.500 3613.980 1143.740 ;
  LAYER metal2 ;
  RECT 3612.860 1140.500 3613.980 1143.740 ;
  LAYER metal1 ;
  RECT 3612.860 1140.500 3613.980 1143.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1132.660 3613.980 1135.900 ;
  LAYER metal4 ;
  RECT 3612.860 1132.660 3613.980 1135.900 ;
  LAYER metal3 ;
  RECT 3612.860 1132.660 3613.980 1135.900 ;
  LAYER metal2 ;
  RECT 3612.860 1132.660 3613.980 1135.900 ;
  LAYER metal1 ;
  RECT 3612.860 1132.660 3613.980 1135.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1124.820 3613.980 1128.060 ;
  LAYER metal4 ;
  RECT 3612.860 1124.820 3613.980 1128.060 ;
  LAYER metal3 ;
  RECT 3612.860 1124.820 3613.980 1128.060 ;
  LAYER metal2 ;
  RECT 3612.860 1124.820 3613.980 1128.060 ;
  LAYER metal1 ;
  RECT 3612.860 1124.820 3613.980 1128.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1116.980 3613.980 1120.220 ;
  LAYER metal4 ;
  RECT 3612.860 1116.980 3613.980 1120.220 ;
  LAYER metal3 ;
  RECT 3612.860 1116.980 3613.980 1120.220 ;
  LAYER metal2 ;
  RECT 3612.860 1116.980 3613.980 1120.220 ;
  LAYER metal1 ;
  RECT 3612.860 1116.980 3613.980 1120.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1109.140 3613.980 1112.380 ;
  LAYER metal4 ;
  RECT 3612.860 1109.140 3613.980 1112.380 ;
  LAYER metal3 ;
  RECT 3612.860 1109.140 3613.980 1112.380 ;
  LAYER metal2 ;
  RECT 3612.860 1109.140 3613.980 1112.380 ;
  LAYER metal1 ;
  RECT 3612.860 1109.140 3613.980 1112.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1069.940 3613.980 1073.180 ;
  LAYER metal4 ;
  RECT 3612.860 1069.940 3613.980 1073.180 ;
  LAYER metal3 ;
  RECT 3612.860 1069.940 3613.980 1073.180 ;
  LAYER metal2 ;
  RECT 3612.860 1069.940 3613.980 1073.180 ;
  LAYER metal1 ;
  RECT 3612.860 1069.940 3613.980 1073.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1062.100 3613.980 1065.340 ;
  LAYER metal4 ;
  RECT 3612.860 1062.100 3613.980 1065.340 ;
  LAYER metal3 ;
  RECT 3612.860 1062.100 3613.980 1065.340 ;
  LAYER metal2 ;
  RECT 3612.860 1062.100 3613.980 1065.340 ;
  LAYER metal1 ;
  RECT 3612.860 1062.100 3613.980 1065.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1054.260 3613.980 1057.500 ;
  LAYER metal4 ;
  RECT 3612.860 1054.260 3613.980 1057.500 ;
  LAYER metal3 ;
  RECT 3612.860 1054.260 3613.980 1057.500 ;
  LAYER metal2 ;
  RECT 3612.860 1054.260 3613.980 1057.500 ;
  LAYER metal1 ;
  RECT 3612.860 1054.260 3613.980 1057.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1046.420 3613.980 1049.660 ;
  LAYER metal4 ;
  RECT 3612.860 1046.420 3613.980 1049.660 ;
  LAYER metal3 ;
  RECT 3612.860 1046.420 3613.980 1049.660 ;
  LAYER metal2 ;
  RECT 3612.860 1046.420 3613.980 1049.660 ;
  LAYER metal1 ;
  RECT 3612.860 1046.420 3613.980 1049.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1038.580 3613.980 1041.820 ;
  LAYER metal4 ;
  RECT 3612.860 1038.580 3613.980 1041.820 ;
  LAYER metal3 ;
  RECT 3612.860 1038.580 3613.980 1041.820 ;
  LAYER metal2 ;
  RECT 3612.860 1038.580 3613.980 1041.820 ;
  LAYER metal1 ;
  RECT 3612.860 1038.580 3613.980 1041.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1030.740 3613.980 1033.980 ;
  LAYER metal4 ;
  RECT 3612.860 1030.740 3613.980 1033.980 ;
  LAYER metal3 ;
  RECT 3612.860 1030.740 3613.980 1033.980 ;
  LAYER metal2 ;
  RECT 3612.860 1030.740 3613.980 1033.980 ;
  LAYER metal1 ;
  RECT 3612.860 1030.740 3613.980 1033.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 991.540 3613.980 994.780 ;
  LAYER metal4 ;
  RECT 3612.860 991.540 3613.980 994.780 ;
  LAYER metal3 ;
  RECT 3612.860 991.540 3613.980 994.780 ;
  LAYER metal2 ;
  RECT 3612.860 991.540 3613.980 994.780 ;
  LAYER metal1 ;
  RECT 3612.860 991.540 3613.980 994.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 983.700 3613.980 986.940 ;
  LAYER metal4 ;
  RECT 3612.860 983.700 3613.980 986.940 ;
  LAYER metal3 ;
  RECT 3612.860 983.700 3613.980 986.940 ;
  LAYER metal2 ;
  RECT 3612.860 983.700 3613.980 986.940 ;
  LAYER metal1 ;
  RECT 3612.860 983.700 3613.980 986.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 975.860 3613.980 979.100 ;
  LAYER metal4 ;
  RECT 3612.860 975.860 3613.980 979.100 ;
  LAYER metal3 ;
  RECT 3612.860 975.860 3613.980 979.100 ;
  LAYER metal2 ;
  RECT 3612.860 975.860 3613.980 979.100 ;
  LAYER metal1 ;
  RECT 3612.860 975.860 3613.980 979.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 968.020 3613.980 971.260 ;
  LAYER metal4 ;
  RECT 3612.860 968.020 3613.980 971.260 ;
  LAYER metal3 ;
  RECT 3612.860 968.020 3613.980 971.260 ;
  LAYER metal2 ;
  RECT 3612.860 968.020 3613.980 971.260 ;
  LAYER metal1 ;
  RECT 3612.860 968.020 3613.980 971.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 960.180 3613.980 963.420 ;
  LAYER metal4 ;
  RECT 3612.860 960.180 3613.980 963.420 ;
  LAYER metal3 ;
  RECT 3612.860 960.180 3613.980 963.420 ;
  LAYER metal2 ;
  RECT 3612.860 960.180 3613.980 963.420 ;
  LAYER metal1 ;
  RECT 3612.860 960.180 3613.980 963.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 952.340 3613.980 955.580 ;
  LAYER metal4 ;
  RECT 3612.860 952.340 3613.980 955.580 ;
  LAYER metal3 ;
  RECT 3612.860 952.340 3613.980 955.580 ;
  LAYER metal2 ;
  RECT 3612.860 952.340 3613.980 955.580 ;
  LAYER metal1 ;
  RECT 3612.860 952.340 3613.980 955.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 913.140 3613.980 916.380 ;
  LAYER metal4 ;
  RECT 3612.860 913.140 3613.980 916.380 ;
  LAYER metal3 ;
  RECT 3612.860 913.140 3613.980 916.380 ;
  LAYER metal2 ;
  RECT 3612.860 913.140 3613.980 916.380 ;
  LAYER metal1 ;
  RECT 3612.860 913.140 3613.980 916.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 905.300 3613.980 908.540 ;
  LAYER metal4 ;
  RECT 3612.860 905.300 3613.980 908.540 ;
  LAYER metal3 ;
  RECT 3612.860 905.300 3613.980 908.540 ;
  LAYER metal2 ;
  RECT 3612.860 905.300 3613.980 908.540 ;
  LAYER metal1 ;
  RECT 3612.860 905.300 3613.980 908.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 897.460 3613.980 900.700 ;
  LAYER metal4 ;
  RECT 3612.860 897.460 3613.980 900.700 ;
  LAYER metal3 ;
  RECT 3612.860 897.460 3613.980 900.700 ;
  LAYER metal2 ;
  RECT 3612.860 897.460 3613.980 900.700 ;
  LAYER metal1 ;
  RECT 3612.860 897.460 3613.980 900.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 889.620 3613.980 892.860 ;
  LAYER metal4 ;
  RECT 3612.860 889.620 3613.980 892.860 ;
  LAYER metal3 ;
  RECT 3612.860 889.620 3613.980 892.860 ;
  LAYER metal2 ;
  RECT 3612.860 889.620 3613.980 892.860 ;
  LAYER metal1 ;
  RECT 3612.860 889.620 3613.980 892.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 881.780 3613.980 885.020 ;
  LAYER metal4 ;
  RECT 3612.860 881.780 3613.980 885.020 ;
  LAYER metal3 ;
  RECT 3612.860 881.780 3613.980 885.020 ;
  LAYER metal2 ;
  RECT 3612.860 881.780 3613.980 885.020 ;
  LAYER metal1 ;
  RECT 3612.860 881.780 3613.980 885.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 873.940 3613.980 877.180 ;
  LAYER metal4 ;
  RECT 3612.860 873.940 3613.980 877.180 ;
  LAYER metal3 ;
  RECT 3612.860 873.940 3613.980 877.180 ;
  LAYER metal2 ;
  RECT 3612.860 873.940 3613.980 877.180 ;
  LAYER metal1 ;
  RECT 3612.860 873.940 3613.980 877.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 834.740 3613.980 837.980 ;
  LAYER metal4 ;
  RECT 3612.860 834.740 3613.980 837.980 ;
  LAYER metal3 ;
  RECT 3612.860 834.740 3613.980 837.980 ;
  LAYER metal2 ;
  RECT 3612.860 834.740 3613.980 837.980 ;
  LAYER metal1 ;
  RECT 3612.860 834.740 3613.980 837.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 826.900 3613.980 830.140 ;
  LAYER metal4 ;
  RECT 3612.860 826.900 3613.980 830.140 ;
  LAYER metal3 ;
  RECT 3612.860 826.900 3613.980 830.140 ;
  LAYER metal2 ;
  RECT 3612.860 826.900 3613.980 830.140 ;
  LAYER metal1 ;
  RECT 3612.860 826.900 3613.980 830.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 819.060 3613.980 822.300 ;
  LAYER metal4 ;
  RECT 3612.860 819.060 3613.980 822.300 ;
  LAYER metal3 ;
  RECT 3612.860 819.060 3613.980 822.300 ;
  LAYER metal2 ;
  RECT 3612.860 819.060 3613.980 822.300 ;
  LAYER metal1 ;
  RECT 3612.860 819.060 3613.980 822.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 811.220 3613.980 814.460 ;
  LAYER metal4 ;
  RECT 3612.860 811.220 3613.980 814.460 ;
  LAYER metal3 ;
  RECT 3612.860 811.220 3613.980 814.460 ;
  LAYER metal2 ;
  RECT 3612.860 811.220 3613.980 814.460 ;
  LAYER metal1 ;
  RECT 3612.860 811.220 3613.980 814.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 803.380 3613.980 806.620 ;
  LAYER metal4 ;
  RECT 3612.860 803.380 3613.980 806.620 ;
  LAYER metal3 ;
  RECT 3612.860 803.380 3613.980 806.620 ;
  LAYER metal2 ;
  RECT 3612.860 803.380 3613.980 806.620 ;
  LAYER metal1 ;
  RECT 3612.860 803.380 3613.980 806.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 795.540 3613.980 798.780 ;
  LAYER metal4 ;
  RECT 3612.860 795.540 3613.980 798.780 ;
  LAYER metal3 ;
  RECT 3612.860 795.540 3613.980 798.780 ;
  LAYER metal2 ;
  RECT 3612.860 795.540 3613.980 798.780 ;
  LAYER metal1 ;
  RECT 3612.860 795.540 3613.980 798.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 756.340 3613.980 759.580 ;
  LAYER metal4 ;
  RECT 3612.860 756.340 3613.980 759.580 ;
  LAYER metal3 ;
  RECT 3612.860 756.340 3613.980 759.580 ;
  LAYER metal2 ;
  RECT 3612.860 756.340 3613.980 759.580 ;
  LAYER metal1 ;
  RECT 3612.860 756.340 3613.980 759.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 748.500 3613.980 751.740 ;
  LAYER metal4 ;
  RECT 3612.860 748.500 3613.980 751.740 ;
  LAYER metal3 ;
  RECT 3612.860 748.500 3613.980 751.740 ;
  LAYER metal2 ;
  RECT 3612.860 748.500 3613.980 751.740 ;
  LAYER metal1 ;
  RECT 3612.860 748.500 3613.980 751.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 740.660 3613.980 743.900 ;
  LAYER metal4 ;
  RECT 3612.860 740.660 3613.980 743.900 ;
  LAYER metal3 ;
  RECT 3612.860 740.660 3613.980 743.900 ;
  LAYER metal2 ;
  RECT 3612.860 740.660 3613.980 743.900 ;
  LAYER metal1 ;
  RECT 3612.860 740.660 3613.980 743.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 732.820 3613.980 736.060 ;
  LAYER metal4 ;
  RECT 3612.860 732.820 3613.980 736.060 ;
  LAYER metal3 ;
  RECT 3612.860 732.820 3613.980 736.060 ;
  LAYER metal2 ;
  RECT 3612.860 732.820 3613.980 736.060 ;
  LAYER metal1 ;
  RECT 3612.860 732.820 3613.980 736.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 724.980 3613.980 728.220 ;
  LAYER metal4 ;
  RECT 3612.860 724.980 3613.980 728.220 ;
  LAYER metal3 ;
  RECT 3612.860 724.980 3613.980 728.220 ;
  LAYER metal2 ;
  RECT 3612.860 724.980 3613.980 728.220 ;
  LAYER metal1 ;
  RECT 3612.860 724.980 3613.980 728.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 717.140 3613.980 720.380 ;
  LAYER metal4 ;
  RECT 3612.860 717.140 3613.980 720.380 ;
  LAYER metal3 ;
  RECT 3612.860 717.140 3613.980 720.380 ;
  LAYER metal2 ;
  RECT 3612.860 717.140 3613.980 720.380 ;
  LAYER metal1 ;
  RECT 3612.860 717.140 3613.980 720.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 677.940 3613.980 681.180 ;
  LAYER metal4 ;
  RECT 3612.860 677.940 3613.980 681.180 ;
  LAYER metal3 ;
  RECT 3612.860 677.940 3613.980 681.180 ;
  LAYER metal2 ;
  RECT 3612.860 677.940 3613.980 681.180 ;
  LAYER metal1 ;
  RECT 3612.860 677.940 3613.980 681.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 670.100 3613.980 673.340 ;
  LAYER metal4 ;
  RECT 3612.860 670.100 3613.980 673.340 ;
  LAYER metal3 ;
  RECT 3612.860 670.100 3613.980 673.340 ;
  LAYER metal2 ;
  RECT 3612.860 670.100 3613.980 673.340 ;
  LAYER metal1 ;
  RECT 3612.860 670.100 3613.980 673.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 662.260 3613.980 665.500 ;
  LAYER metal4 ;
  RECT 3612.860 662.260 3613.980 665.500 ;
  LAYER metal3 ;
  RECT 3612.860 662.260 3613.980 665.500 ;
  LAYER metal2 ;
  RECT 3612.860 662.260 3613.980 665.500 ;
  LAYER metal1 ;
  RECT 3612.860 662.260 3613.980 665.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 654.420 3613.980 657.660 ;
  LAYER metal4 ;
  RECT 3612.860 654.420 3613.980 657.660 ;
  LAYER metal3 ;
  RECT 3612.860 654.420 3613.980 657.660 ;
  LAYER metal2 ;
  RECT 3612.860 654.420 3613.980 657.660 ;
  LAYER metal1 ;
  RECT 3612.860 654.420 3613.980 657.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 646.580 3613.980 649.820 ;
  LAYER metal4 ;
  RECT 3612.860 646.580 3613.980 649.820 ;
  LAYER metal3 ;
  RECT 3612.860 646.580 3613.980 649.820 ;
  LAYER metal2 ;
  RECT 3612.860 646.580 3613.980 649.820 ;
  LAYER metal1 ;
  RECT 3612.860 646.580 3613.980 649.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 638.740 3613.980 641.980 ;
  LAYER metal4 ;
  RECT 3612.860 638.740 3613.980 641.980 ;
  LAYER metal3 ;
  RECT 3612.860 638.740 3613.980 641.980 ;
  LAYER metal2 ;
  RECT 3612.860 638.740 3613.980 641.980 ;
  LAYER metal1 ;
  RECT 3612.860 638.740 3613.980 641.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 599.540 3613.980 602.780 ;
  LAYER metal4 ;
  RECT 3612.860 599.540 3613.980 602.780 ;
  LAYER metal3 ;
  RECT 3612.860 599.540 3613.980 602.780 ;
  LAYER metal2 ;
  RECT 3612.860 599.540 3613.980 602.780 ;
  LAYER metal1 ;
  RECT 3612.860 599.540 3613.980 602.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 591.700 3613.980 594.940 ;
  LAYER metal4 ;
  RECT 3612.860 591.700 3613.980 594.940 ;
  LAYER metal3 ;
  RECT 3612.860 591.700 3613.980 594.940 ;
  LAYER metal2 ;
  RECT 3612.860 591.700 3613.980 594.940 ;
  LAYER metal1 ;
  RECT 3612.860 591.700 3613.980 594.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 583.860 3613.980 587.100 ;
  LAYER metal4 ;
  RECT 3612.860 583.860 3613.980 587.100 ;
  LAYER metal3 ;
  RECT 3612.860 583.860 3613.980 587.100 ;
  LAYER metal2 ;
  RECT 3612.860 583.860 3613.980 587.100 ;
  LAYER metal1 ;
  RECT 3612.860 583.860 3613.980 587.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 576.020 3613.980 579.260 ;
  LAYER metal4 ;
  RECT 3612.860 576.020 3613.980 579.260 ;
  LAYER metal3 ;
  RECT 3612.860 576.020 3613.980 579.260 ;
  LAYER metal2 ;
  RECT 3612.860 576.020 3613.980 579.260 ;
  LAYER metal1 ;
  RECT 3612.860 576.020 3613.980 579.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 568.180 3613.980 571.420 ;
  LAYER metal4 ;
  RECT 3612.860 568.180 3613.980 571.420 ;
  LAYER metal3 ;
  RECT 3612.860 568.180 3613.980 571.420 ;
  LAYER metal2 ;
  RECT 3612.860 568.180 3613.980 571.420 ;
  LAYER metal1 ;
  RECT 3612.860 568.180 3613.980 571.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 560.340 3613.980 563.580 ;
  LAYER metal4 ;
  RECT 3612.860 560.340 3613.980 563.580 ;
  LAYER metal3 ;
  RECT 3612.860 560.340 3613.980 563.580 ;
  LAYER metal2 ;
  RECT 3612.860 560.340 3613.980 563.580 ;
  LAYER metal1 ;
  RECT 3612.860 560.340 3613.980 563.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 521.140 3613.980 524.380 ;
  LAYER metal4 ;
  RECT 3612.860 521.140 3613.980 524.380 ;
  LAYER metal3 ;
  RECT 3612.860 521.140 3613.980 524.380 ;
  LAYER metal2 ;
  RECT 3612.860 521.140 3613.980 524.380 ;
  LAYER metal1 ;
  RECT 3612.860 521.140 3613.980 524.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 513.300 3613.980 516.540 ;
  LAYER metal4 ;
  RECT 3612.860 513.300 3613.980 516.540 ;
  LAYER metal3 ;
  RECT 3612.860 513.300 3613.980 516.540 ;
  LAYER metal2 ;
  RECT 3612.860 513.300 3613.980 516.540 ;
  LAYER metal1 ;
  RECT 3612.860 513.300 3613.980 516.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 505.460 3613.980 508.700 ;
  LAYER metal4 ;
  RECT 3612.860 505.460 3613.980 508.700 ;
  LAYER metal3 ;
  RECT 3612.860 505.460 3613.980 508.700 ;
  LAYER metal2 ;
  RECT 3612.860 505.460 3613.980 508.700 ;
  LAYER metal1 ;
  RECT 3612.860 505.460 3613.980 508.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 497.620 3613.980 500.860 ;
  LAYER metal4 ;
  RECT 3612.860 497.620 3613.980 500.860 ;
  LAYER metal3 ;
  RECT 3612.860 497.620 3613.980 500.860 ;
  LAYER metal2 ;
  RECT 3612.860 497.620 3613.980 500.860 ;
  LAYER metal1 ;
  RECT 3612.860 497.620 3613.980 500.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 489.780 3613.980 493.020 ;
  LAYER metal4 ;
  RECT 3612.860 489.780 3613.980 493.020 ;
  LAYER metal3 ;
  RECT 3612.860 489.780 3613.980 493.020 ;
  LAYER metal2 ;
  RECT 3612.860 489.780 3613.980 493.020 ;
  LAYER metal1 ;
  RECT 3612.860 489.780 3613.980 493.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 481.940 3613.980 485.180 ;
  LAYER metal4 ;
  RECT 3612.860 481.940 3613.980 485.180 ;
  LAYER metal3 ;
  RECT 3612.860 481.940 3613.980 485.180 ;
  LAYER metal2 ;
  RECT 3612.860 481.940 3613.980 485.180 ;
  LAYER metal1 ;
  RECT 3612.860 481.940 3613.980 485.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 442.740 3613.980 445.980 ;
  LAYER metal4 ;
  RECT 3612.860 442.740 3613.980 445.980 ;
  LAYER metal3 ;
  RECT 3612.860 442.740 3613.980 445.980 ;
  LAYER metal2 ;
  RECT 3612.860 442.740 3613.980 445.980 ;
  LAYER metal1 ;
  RECT 3612.860 442.740 3613.980 445.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 434.900 3613.980 438.140 ;
  LAYER metal4 ;
  RECT 3612.860 434.900 3613.980 438.140 ;
  LAYER metal3 ;
  RECT 3612.860 434.900 3613.980 438.140 ;
  LAYER metal2 ;
  RECT 3612.860 434.900 3613.980 438.140 ;
  LAYER metal1 ;
  RECT 3612.860 434.900 3613.980 438.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 427.060 3613.980 430.300 ;
  LAYER metal4 ;
  RECT 3612.860 427.060 3613.980 430.300 ;
  LAYER metal3 ;
  RECT 3612.860 427.060 3613.980 430.300 ;
  LAYER metal2 ;
  RECT 3612.860 427.060 3613.980 430.300 ;
  LAYER metal1 ;
  RECT 3612.860 427.060 3613.980 430.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 419.220 3613.980 422.460 ;
  LAYER metal4 ;
  RECT 3612.860 419.220 3613.980 422.460 ;
  LAYER metal3 ;
  RECT 3612.860 419.220 3613.980 422.460 ;
  LAYER metal2 ;
  RECT 3612.860 419.220 3613.980 422.460 ;
  LAYER metal1 ;
  RECT 3612.860 419.220 3613.980 422.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 411.380 3613.980 414.620 ;
  LAYER metal4 ;
  RECT 3612.860 411.380 3613.980 414.620 ;
  LAYER metal3 ;
  RECT 3612.860 411.380 3613.980 414.620 ;
  LAYER metal2 ;
  RECT 3612.860 411.380 3613.980 414.620 ;
  LAYER metal1 ;
  RECT 3612.860 411.380 3613.980 414.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 403.540 3613.980 406.780 ;
  LAYER metal4 ;
  RECT 3612.860 403.540 3613.980 406.780 ;
  LAYER metal3 ;
  RECT 3612.860 403.540 3613.980 406.780 ;
  LAYER metal2 ;
  RECT 3612.860 403.540 3613.980 406.780 ;
  LAYER metal1 ;
  RECT 3612.860 403.540 3613.980 406.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 364.340 3613.980 367.580 ;
  LAYER metal4 ;
  RECT 3612.860 364.340 3613.980 367.580 ;
  LAYER metal3 ;
  RECT 3612.860 364.340 3613.980 367.580 ;
  LAYER metal2 ;
  RECT 3612.860 364.340 3613.980 367.580 ;
  LAYER metal1 ;
  RECT 3612.860 364.340 3613.980 367.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 356.500 3613.980 359.740 ;
  LAYER metal4 ;
  RECT 3612.860 356.500 3613.980 359.740 ;
  LAYER metal3 ;
  RECT 3612.860 356.500 3613.980 359.740 ;
  LAYER metal2 ;
  RECT 3612.860 356.500 3613.980 359.740 ;
  LAYER metal1 ;
  RECT 3612.860 356.500 3613.980 359.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 348.660 3613.980 351.900 ;
  LAYER metal4 ;
  RECT 3612.860 348.660 3613.980 351.900 ;
  LAYER metal3 ;
  RECT 3612.860 348.660 3613.980 351.900 ;
  LAYER metal2 ;
  RECT 3612.860 348.660 3613.980 351.900 ;
  LAYER metal1 ;
  RECT 3612.860 348.660 3613.980 351.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 340.820 3613.980 344.060 ;
  LAYER metal4 ;
  RECT 3612.860 340.820 3613.980 344.060 ;
  LAYER metal3 ;
  RECT 3612.860 340.820 3613.980 344.060 ;
  LAYER metal2 ;
  RECT 3612.860 340.820 3613.980 344.060 ;
  LAYER metal1 ;
  RECT 3612.860 340.820 3613.980 344.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 332.980 3613.980 336.220 ;
  LAYER metal4 ;
  RECT 3612.860 332.980 3613.980 336.220 ;
  LAYER metal3 ;
  RECT 3612.860 332.980 3613.980 336.220 ;
  LAYER metal2 ;
  RECT 3612.860 332.980 3613.980 336.220 ;
  LAYER metal1 ;
  RECT 3612.860 332.980 3613.980 336.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 325.140 3613.980 328.380 ;
  LAYER metal4 ;
  RECT 3612.860 325.140 3613.980 328.380 ;
  LAYER metal3 ;
  RECT 3612.860 325.140 3613.980 328.380 ;
  LAYER metal2 ;
  RECT 3612.860 325.140 3613.980 328.380 ;
  LAYER metal1 ;
  RECT 3612.860 325.140 3613.980 328.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 285.940 3613.980 289.180 ;
  LAYER metal4 ;
  RECT 3612.860 285.940 3613.980 289.180 ;
  LAYER metal3 ;
  RECT 3612.860 285.940 3613.980 289.180 ;
  LAYER metal2 ;
  RECT 3612.860 285.940 3613.980 289.180 ;
  LAYER metal1 ;
  RECT 3612.860 285.940 3613.980 289.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 278.100 3613.980 281.340 ;
  LAYER metal4 ;
  RECT 3612.860 278.100 3613.980 281.340 ;
  LAYER metal3 ;
  RECT 3612.860 278.100 3613.980 281.340 ;
  LAYER metal2 ;
  RECT 3612.860 278.100 3613.980 281.340 ;
  LAYER metal1 ;
  RECT 3612.860 278.100 3613.980 281.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 270.260 3613.980 273.500 ;
  LAYER metal4 ;
  RECT 3612.860 270.260 3613.980 273.500 ;
  LAYER metal3 ;
  RECT 3612.860 270.260 3613.980 273.500 ;
  LAYER metal2 ;
  RECT 3612.860 270.260 3613.980 273.500 ;
  LAYER metal1 ;
  RECT 3612.860 270.260 3613.980 273.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 262.420 3613.980 265.660 ;
  LAYER metal4 ;
  RECT 3612.860 262.420 3613.980 265.660 ;
  LAYER metal3 ;
  RECT 3612.860 262.420 3613.980 265.660 ;
  LAYER metal2 ;
  RECT 3612.860 262.420 3613.980 265.660 ;
  LAYER metal1 ;
  RECT 3612.860 262.420 3613.980 265.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 254.580 3613.980 257.820 ;
  LAYER metal4 ;
  RECT 3612.860 254.580 3613.980 257.820 ;
  LAYER metal3 ;
  RECT 3612.860 254.580 3613.980 257.820 ;
  LAYER metal2 ;
  RECT 3612.860 254.580 3613.980 257.820 ;
  LAYER metal1 ;
  RECT 3612.860 254.580 3613.980 257.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 246.740 3613.980 249.980 ;
  LAYER metal4 ;
  RECT 3612.860 246.740 3613.980 249.980 ;
  LAYER metal3 ;
  RECT 3612.860 246.740 3613.980 249.980 ;
  LAYER metal2 ;
  RECT 3612.860 246.740 3613.980 249.980 ;
  LAYER metal1 ;
  RECT 3612.860 246.740 3613.980 249.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 207.540 3613.980 210.780 ;
  LAYER metal4 ;
  RECT 3612.860 207.540 3613.980 210.780 ;
  LAYER metal3 ;
  RECT 3612.860 207.540 3613.980 210.780 ;
  LAYER metal2 ;
  RECT 3612.860 207.540 3613.980 210.780 ;
  LAYER metal1 ;
  RECT 3612.860 207.540 3613.980 210.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 199.700 3613.980 202.940 ;
  LAYER metal4 ;
  RECT 3612.860 199.700 3613.980 202.940 ;
  LAYER metal3 ;
  RECT 3612.860 199.700 3613.980 202.940 ;
  LAYER metal2 ;
  RECT 3612.860 199.700 3613.980 202.940 ;
  LAYER metal1 ;
  RECT 3612.860 199.700 3613.980 202.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 191.860 3613.980 195.100 ;
  LAYER metal4 ;
  RECT 3612.860 191.860 3613.980 195.100 ;
  LAYER metal3 ;
  RECT 3612.860 191.860 3613.980 195.100 ;
  LAYER metal2 ;
  RECT 3612.860 191.860 3613.980 195.100 ;
  LAYER metal1 ;
  RECT 3612.860 191.860 3613.980 195.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 184.020 3613.980 187.260 ;
  LAYER metal4 ;
  RECT 3612.860 184.020 3613.980 187.260 ;
  LAYER metal3 ;
  RECT 3612.860 184.020 3613.980 187.260 ;
  LAYER metal2 ;
  RECT 3612.860 184.020 3613.980 187.260 ;
  LAYER metal1 ;
  RECT 3612.860 184.020 3613.980 187.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 176.180 3613.980 179.420 ;
  LAYER metal4 ;
  RECT 3612.860 176.180 3613.980 179.420 ;
  LAYER metal3 ;
  RECT 3612.860 176.180 3613.980 179.420 ;
  LAYER metal2 ;
  RECT 3612.860 176.180 3613.980 179.420 ;
  LAYER metal1 ;
  RECT 3612.860 176.180 3613.980 179.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 168.340 3613.980 171.580 ;
  LAYER metal4 ;
  RECT 3612.860 168.340 3613.980 171.580 ;
  LAYER metal3 ;
  RECT 3612.860 168.340 3613.980 171.580 ;
  LAYER metal2 ;
  RECT 3612.860 168.340 3613.980 171.580 ;
  LAYER metal1 ;
  RECT 3612.860 168.340 3613.980 171.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 129.140 3613.980 132.380 ;
  LAYER metal4 ;
  RECT 3612.860 129.140 3613.980 132.380 ;
  LAYER metal3 ;
  RECT 3612.860 129.140 3613.980 132.380 ;
  LAYER metal2 ;
  RECT 3612.860 129.140 3613.980 132.380 ;
  LAYER metal1 ;
  RECT 3612.860 129.140 3613.980 132.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 121.300 3613.980 124.540 ;
  LAYER metal4 ;
  RECT 3612.860 121.300 3613.980 124.540 ;
  LAYER metal3 ;
  RECT 3612.860 121.300 3613.980 124.540 ;
  LAYER metal2 ;
  RECT 3612.860 121.300 3613.980 124.540 ;
  LAYER metal1 ;
  RECT 3612.860 121.300 3613.980 124.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 113.460 3613.980 116.700 ;
  LAYER metal4 ;
  RECT 3612.860 113.460 3613.980 116.700 ;
  LAYER metal3 ;
  RECT 3612.860 113.460 3613.980 116.700 ;
  LAYER metal2 ;
  RECT 3612.860 113.460 3613.980 116.700 ;
  LAYER metal1 ;
  RECT 3612.860 113.460 3613.980 116.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 105.620 3613.980 108.860 ;
  LAYER metal4 ;
  RECT 3612.860 105.620 3613.980 108.860 ;
  LAYER metal3 ;
  RECT 3612.860 105.620 3613.980 108.860 ;
  LAYER metal2 ;
  RECT 3612.860 105.620 3613.980 108.860 ;
  LAYER metal1 ;
  RECT 3612.860 105.620 3613.980 108.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 97.780 3613.980 101.020 ;
  LAYER metal4 ;
  RECT 3612.860 97.780 3613.980 101.020 ;
  LAYER metal3 ;
  RECT 3612.860 97.780 3613.980 101.020 ;
  LAYER metal2 ;
  RECT 3612.860 97.780 3613.980 101.020 ;
  LAYER metal1 ;
  RECT 3612.860 97.780 3613.980 101.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 89.940 3613.980 93.180 ;
  LAYER metal4 ;
  RECT 3612.860 89.940 3613.980 93.180 ;
  LAYER metal3 ;
  RECT 3612.860 89.940 3613.980 93.180 ;
  LAYER metal2 ;
  RECT 3612.860 89.940 3613.980 93.180 ;
  LAYER metal1 ;
  RECT 3612.860 89.940 3613.980 93.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 50.740 3613.980 53.980 ;
  LAYER metal4 ;
  RECT 3612.860 50.740 3613.980 53.980 ;
  LAYER metal3 ;
  RECT 3612.860 50.740 3613.980 53.980 ;
  LAYER metal2 ;
  RECT 3612.860 50.740 3613.980 53.980 ;
  LAYER metal1 ;
  RECT 3612.860 50.740 3613.980 53.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 42.900 3613.980 46.140 ;
  LAYER metal4 ;
  RECT 3612.860 42.900 3613.980 46.140 ;
  LAYER metal3 ;
  RECT 3612.860 42.900 3613.980 46.140 ;
  LAYER metal2 ;
  RECT 3612.860 42.900 3613.980 46.140 ;
  LAYER metal1 ;
  RECT 3612.860 42.900 3613.980 46.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 35.060 3613.980 38.300 ;
  LAYER metal4 ;
  RECT 3612.860 35.060 3613.980 38.300 ;
  LAYER metal3 ;
  RECT 3612.860 35.060 3613.980 38.300 ;
  LAYER metal2 ;
  RECT 3612.860 35.060 3613.980 38.300 ;
  LAYER metal1 ;
  RECT 3612.860 35.060 3613.980 38.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 27.220 3613.980 30.460 ;
  LAYER metal4 ;
  RECT 3612.860 27.220 3613.980 30.460 ;
  LAYER metal3 ;
  RECT 3612.860 27.220 3613.980 30.460 ;
  LAYER metal2 ;
  RECT 3612.860 27.220 3613.980 30.460 ;
  LAYER metal1 ;
  RECT 3612.860 27.220 3613.980 30.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 19.380 3613.980 22.620 ;
  LAYER metal4 ;
  RECT 3612.860 19.380 3613.980 22.620 ;
  LAYER metal3 ;
  RECT 3612.860 19.380 3613.980 22.620 ;
  LAYER metal2 ;
  RECT 3612.860 19.380 3613.980 22.620 ;
  LAYER metal1 ;
  RECT 3612.860 19.380 3613.980 22.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 11.540 3613.980 14.780 ;
  LAYER metal4 ;
  RECT 3612.860 11.540 3613.980 14.780 ;
  LAYER metal3 ;
  RECT 3612.860 11.540 3613.980 14.780 ;
  LAYER metal2 ;
  RECT 3612.860 11.540 3613.980 14.780 ;
  LAYER metal1 ;
  RECT 3612.860 11.540 3613.980 14.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1697.140 1.120 1700.380 ;
  LAYER metal4 ;
  RECT 0.000 1697.140 1.120 1700.380 ;
  LAYER metal3 ;
  RECT 0.000 1697.140 1.120 1700.380 ;
  LAYER metal2 ;
  RECT 0.000 1697.140 1.120 1700.380 ;
  LAYER metal1 ;
  RECT 0.000 1697.140 1.120 1700.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1689.300 1.120 1692.540 ;
  LAYER metal4 ;
  RECT 0.000 1689.300 1.120 1692.540 ;
  LAYER metal3 ;
  RECT 0.000 1689.300 1.120 1692.540 ;
  LAYER metal2 ;
  RECT 0.000 1689.300 1.120 1692.540 ;
  LAYER metal1 ;
  RECT 0.000 1689.300 1.120 1692.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1681.460 1.120 1684.700 ;
  LAYER metal4 ;
  RECT 0.000 1681.460 1.120 1684.700 ;
  LAYER metal3 ;
  RECT 0.000 1681.460 1.120 1684.700 ;
  LAYER metal2 ;
  RECT 0.000 1681.460 1.120 1684.700 ;
  LAYER metal1 ;
  RECT 0.000 1681.460 1.120 1684.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1673.620 1.120 1676.860 ;
  LAYER metal4 ;
  RECT 0.000 1673.620 1.120 1676.860 ;
  LAYER metal3 ;
  RECT 0.000 1673.620 1.120 1676.860 ;
  LAYER metal2 ;
  RECT 0.000 1673.620 1.120 1676.860 ;
  LAYER metal1 ;
  RECT 0.000 1673.620 1.120 1676.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1665.780 1.120 1669.020 ;
  LAYER metal4 ;
  RECT 0.000 1665.780 1.120 1669.020 ;
  LAYER metal3 ;
  RECT 0.000 1665.780 1.120 1669.020 ;
  LAYER metal2 ;
  RECT 0.000 1665.780 1.120 1669.020 ;
  LAYER metal1 ;
  RECT 0.000 1665.780 1.120 1669.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1657.940 1.120 1661.180 ;
  LAYER metal4 ;
  RECT 0.000 1657.940 1.120 1661.180 ;
  LAYER metal3 ;
  RECT 0.000 1657.940 1.120 1661.180 ;
  LAYER metal2 ;
  RECT 0.000 1657.940 1.120 1661.180 ;
  LAYER metal1 ;
  RECT 0.000 1657.940 1.120 1661.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1618.740 1.120 1621.980 ;
  LAYER metal4 ;
  RECT 0.000 1618.740 1.120 1621.980 ;
  LAYER metal3 ;
  RECT 0.000 1618.740 1.120 1621.980 ;
  LAYER metal2 ;
  RECT 0.000 1618.740 1.120 1621.980 ;
  LAYER metal1 ;
  RECT 0.000 1618.740 1.120 1621.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1610.900 1.120 1614.140 ;
  LAYER metal4 ;
  RECT 0.000 1610.900 1.120 1614.140 ;
  LAYER metal3 ;
  RECT 0.000 1610.900 1.120 1614.140 ;
  LAYER metal2 ;
  RECT 0.000 1610.900 1.120 1614.140 ;
  LAYER metal1 ;
  RECT 0.000 1610.900 1.120 1614.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1603.060 1.120 1606.300 ;
  LAYER metal4 ;
  RECT 0.000 1603.060 1.120 1606.300 ;
  LAYER metal3 ;
  RECT 0.000 1603.060 1.120 1606.300 ;
  LAYER metal2 ;
  RECT 0.000 1603.060 1.120 1606.300 ;
  LAYER metal1 ;
  RECT 0.000 1603.060 1.120 1606.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1595.220 1.120 1598.460 ;
  LAYER metal4 ;
  RECT 0.000 1595.220 1.120 1598.460 ;
  LAYER metal3 ;
  RECT 0.000 1595.220 1.120 1598.460 ;
  LAYER metal2 ;
  RECT 0.000 1595.220 1.120 1598.460 ;
  LAYER metal1 ;
  RECT 0.000 1595.220 1.120 1598.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1587.380 1.120 1590.620 ;
  LAYER metal4 ;
  RECT 0.000 1587.380 1.120 1590.620 ;
  LAYER metal3 ;
  RECT 0.000 1587.380 1.120 1590.620 ;
  LAYER metal2 ;
  RECT 0.000 1587.380 1.120 1590.620 ;
  LAYER metal1 ;
  RECT 0.000 1587.380 1.120 1590.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1579.540 1.120 1582.780 ;
  LAYER metal4 ;
  RECT 0.000 1579.540 1.120 1582.780 ;
  LAYER metal3 ;
  RECT 0.000 1579.540 1.120 1582.780 ;
  LAYER metal2 ;
  RECT 0.000 1579.540 1.120 1582.780 ;
  LAYER metal1 ;
  RECT 0.000 1579.540 1.120 1582.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1540.340 1.120 1543.580 ;
  LAYER metal4 ;
  RECT 0.000 1540.340 1.120 1543.580 ;
  LAYER metal3 ;
  RECT 0.000 1540.340 1.120 1543.580 ;
  LAYER metal2 ;
  RECT 0.000 1540.340 1.120 1543.580 ;
  LAYER metal1 ;
  RECT 0.000 1540.340 1.120 1543.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1532.500 1.120 1535.740 ;
  LAYER metal4 ;
  RECT 0.000 1532.500 1.120 1535.740 ;
  LAYER metal3 ;
  RECT 0.000 1532.500 1.120 1535.740 ;
  LAYER metal2 ;
  RECT 0.000 1532.500 1.120 1535.740 ;
  LAYER metal1 ;
  RECT 0.000 1532.500 1.120 1535.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1524.660 1.120 1527.900 ;
  LAYER metal4 ;
  RECT 0.000 1524.660 1.120 1527.900 ;
  LAYER metal3 ;
  RECT 0.000 1524.660 1.120 1527.900 ;
  LAYER metal2 ;
  RECT 0.000 1524.660 1.120 1527.900 ;
  LAYER metal1 ;
  RECT 0.000 1524.660 1.120 1527.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1516.820 1.120 1520.060 ;
  LAYER metal4 ;
  RECT 0.000 1516.820 1.120 1520.060 ;
  LAYER metal3 ;
  RECT 0.000 1516.820 1.120 1520.060 ;
  LAYER metal2 ;
  RECT 0.000 1516.820 1.120 1520.060 ;
  LAYER metal1 ;
  RECT 0.000 1516.820 1.120 1520.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1508.980 1.120 1512.220 ;
  LAYER metal4 ;
  RECT 0.000 1508.980 1.120 1512.220 ;
  LAYER metal3 ;
  RECT 0.000 1508.980 1.120 1512.220 ;
  LAYER metal2 ;
  RECT 0.000 1508.980 1.120 1512.220 ;
  LAYER metal1 ;
  RECT 0.000 1508.980 1.120 1512.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1501.140 1.120 1504.380 ;
  LAYER metal4 ;
  RECT 0.000 1501.140 1.120 1504.380 ;
  LAYER metal3 ;
  RECT 0.000 1501.140 1.120 1504.380 ;
  LAYER metal2 ;
  RECT 0.000 1501.140 1.120 1504.380 ;
  LAYER metal1 ;
  RECT 0.000 1501.140 1.120 1504.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1461.940 1.120 1465.180 ;
  LAYER metal4 ;
  RECT 0.000 1461.940 1.120 1465.180 ;
  LAYER metal3 ;
  RECT 0.000 1461.940 1.120 1465.180 ;
  LAYER metal2 ;
  RECT 0.000 1461.940 1.120 1465.180 ;
  LAYER metal1 ;
  RECT 0.000 1461.940 1.120 1465.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1454.100 1.120 1457.340 ;
  LAYER metal4 ;
  RECT 0.000 1454.100 1.120 1457.340 ;
  LAYER metal3 ;
  RECT 0.000 1454.100 1.120 1457.340 ;
  LAYER metal2 ;
  RECT 0.000 1454.100 1.120 1457.340 ;
  LAYER metal1 ;
  RECT 0.000 1454.100 1.120 1457.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1446.260 1.120 1449.500 ;
  LAYER metal4 ;
  RECT 0.000 1446.260 1.120 1449.500 ;
  LAYER metal3 ;
  RECT 0.000 1446.260 1.120 1449.500 ;
  LAYER metal2 ;
  RECT 0.000 1446.260 1.120 1449.500 ;
  LAYER metal1 ;
  RECT 0.000 1446.260 1.120 1449.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1438.420 1.120 1441.660 ;
  LAYER metal4 ;
  RECT 0.000 1438.420 1.120 1441.660 ;
  LAYER metal3 ;
  RECT 0.000 1438.420 1.120 1441.660 ;
  LAYER metal2 ;
  RECT 0.000 1438.420 1.120 1441.660 ;
  LAYER metal1 ;
  RECT 0.000 1438.420 1.120 1441.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1430.580 1.120 1433.820 ;
  LAYER metal4 ;
  RECT 0.000 1430.580 1.120 1433.820 ;
  LAYER metal3 ;
  RECT 0.000 1430.580 1.120 1433.820 ;
  LAYER metal2 ;
  RECT 0.000 1430.580 1.120 1433.820 ;
  LAYER metal1 ;
  RECT 0.000 1430.580 1.120 1433.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1422.740 1.120 1425.980 ;
  LAYER metal4 ;
  RECT 0.000 1422.740 1.120 1425.980 ;
  LAYER metal3 ;
  RECT 0.000 1422.740 1.120 1425.980 ;
  LAYER metal2 ;
  RECT 0.000 1422.740 1.120 1425.980 ;
  LAYER metal1 ;
  RECT 0.000 1422.740 1.120 1425.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1383.540 1.120 1386.780 ;
  LAYER metal4 ;
  RECT 0.000 1383.540 1.120 1386.780 ;
  LAYER metal3 ;
  RECT 0.000 1383.540 1.120 1386.780 ;
  LAYER metal2 ;
  RECT 0.000 1383.540 1.120 1386.780 ;
  LAYER metal1 ;
  RECT 0.000 1383.540 1.120 1386.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1375.700 1.120 1378.940 ;
  LAYER metal4 ;
  RECT 0.000 1375.700 1.120 1378.940 ;
  LAYER metal3 ;
  RECT 0.000 1375.700 1.120 1378.940 ;
  LAYER metal2 ;
  RECT 0.000 1375.700 1.120 1378.940 ;
  LAYER metal1 ;
  RECT 0.000 1375.700 1.120 1378.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1367.860 1.120 1371.100 ;
  LAYER metal4 ;
  RECT 0.000 1367.860 1.120 1371.100 ;
  LAYER metal3 ;
  RECT 0.000 1367.860 1.120 1371.100 ;
  LAYER metal2 ;
  RECT 0.000 1367.860 1.120 1371.100 ;
  LAYER metal1 ;
  RECT 0.000 1367.860 1.120 1371.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1360.020 1.120 1363.260 ;
  LAYER metal4 ;
  RECT 0.000 1360.020 1.120 1363.260 ;
  LAYER metal3 ;
  RECT 0.000 1360.020 1.120 1363.260 ;
  LAYER metal2 ;
  RECT 0.000 1360.020 1.120 1363.260 ;
  LAYER metal1 ;
  RECT 0.000 1360.020 1.120 1363.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1352.180 1.120 1355.420 ;
  LAYER metal4 ;
  RECT 0.000 1352.180 1.120 1355.420 ;
  LAYER metal3 ;
  RECT 0.000 1352.180 1.120 1355.420 ;
  LAYER metal2 ;
  RECT 0.000 1352.180 1.120 1355.420 ;
  LAYER metal1 ;
  RECT 0.000 1352.180 1.120 1355.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1344.340 1.120 1347.580 ;
  LAYER metal4 ;
  RECT 0.000 1344.340 1.120 1347.580 ;
  LAYER metal3 ;
  RECT 0.000 1344.340 1.120 1347.580 ;
  LAYER metal2 ;
  RECT 0.000 1344.340 1.120 1347.580 ;
  LAYER metal1 ;
  RECT 0.000 1344.340 1.120 1347.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1305.140 1.120 1308.380 ;
  LAYER metal4 ;
  RECT 0.000 1305.140 1.120 1308.380 ;
  LAYER metal3 ;
  RECT 0.000 1305.140 1.120 1308.380 ;
  LAYER metal2 ;
  RECT 0.000 1305.140 1.120 1308.380 ;
  LAYER metal1 ;
  RECT 0.000 1305.140 1.120 1308.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1297.300 1.120 1300.540 ;
  LAYER metal4 ;
  RECT 0.000 1297.300 1.120 1300.540 ;
  LAYER metal3 ;
  RECT 0.000 1297.300 1.120 1300.540 ;
  LAYER metal2 ;
  RECT 0.000 1297.300 1.120 1300.540 ;
  LAYER metal1 ;
  RECT 0.000 1297.300 1.120 1300.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1289.460 1.120 1292.700 ;
  LAYER metal4 ;
  RECT 0.000 1289.460 1.120 1292.700 ;
  LAYER metal3 ;
  RECT 0.000 1289.460 1.120 1292.700 ;
  LAYER metal2 ;
  RECT 0.000 1289.460 1.120 1292.700 ;
  LAYER metal1 ;
  RECT 0.000 1289.460 1.120 1292.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1281.620 1.120 1284.860 ;
  LAYER metal4 ;
  RECT 0.000 1281.620 1.120 1284.860 ;
  LAYER metal3 ;
  RECT 0.000 1281.620 1.120 1284.860 ;
  LAYER metal2 ;
  RECT 0.000 1281.620 1.120 1284.860 ;
  LAYER metal1 ;
  RECT 0.000 1281.620 1.120 1284.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1273.780 1.120 1277.020 ;
  LAYER metal4 ;
  RECT 0.000 1273.780 1.120 1277.020 ;
  LAYER metal3 ;
  RECT 0.000 1273.780 1.120 1277.020 ;
  LAYER metal2 ;
  RECT 0.000 1273.780 1.120 1277.020 ;
  LAYER metal1 ;
  RECT 0.000 1273.780 1.120 1277.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1265.940 1.120 1269.180 ;
  LAYER metal4 ;
  RECT 0.000 1265.940 1.120 1269.180 ;
  LAYER metal3 ;
  RECT 0.000 1265.940 1.120 1269.180 ;
  LAYER metal2 ;
  RECT 0.000 1265.940 1.120 1269.180 ;
  LAYER metal1 ;
  RECT 0.000 1265.940 1.120 1269.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1226.740 1.120 1229.980 ;
  LAYER metal4 ;
  RECT 0.000 1226.740 1.120 1229.980 ;
  LAYER metal3 ;
  RECT 0.000 1226.740 1.120 1229.980 ;
  LAYER metal2 ;
  RECT 0.000 1226.740 1.120 1229.980 ;
  LAYER metal1 ;
  RECT 0.000 1226.740 1.120 1229.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1218.900 1.120 1222.140 ;
  LAYER metal4 ;
  RECT 0.000 1218.900 1.120 1222.140 ;
  LAYER metal3 ;
  RECT 0.000 1218.900 1.120 1222.140 ;
  LAYER metal2 ;
  RECT 0.000 1218.900 1.120 1222.140 ;
  LAYER metal1 ;
  RECT 0.000 1218.900 1.120 1222.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1211.060 1.120 1214.300 ;
  LAYER metal4 ;
  RECT 0.000 1211.060 1.120 1214.300 ;
  LAYER metal3 ;
  RECT 0.000 1211.060 1.120 1214.300 ;
  LAYER metal2 ;
  RECT 0.000 1211.060 1.120 1214.300 ;
  LAYER metal1 ;
  RECT 0.000 1211.060 1.120 1214.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1203.220 1.120 1206.460 ;
  LAYER metal4 ;
  RECT 0.000 1203.220 1.120 1206.460 ;
  LAYER metal3 ;
  RECT 0.000 1203.220 1.120 1206.460 ;
  LAYER metal2 ;
  RECT 0.000 1203.220 1.120 1206.460 ;
  LAYER metal1 ;
  RECT 0.000 1203.220 1.120 1206.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1195.380 1.120 1198.620 ;
  LAYER metal4 ;
  RECT 0.000 1195.380 1.120 1198.620 ;
  LAYER metal3 ;
  RECT 0.000 1195.380 1.120 1198.620 ;
  LAYER metal2 ;
  RECT 0.000 1195.380 1.120 1198.620 ;
  LAYER metal1 ;
  RECT 0.000 1195.380 1.120 1198.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1187.540 1.120 1190.780 ;
  LAYER metal4 ;
  RECT 0.000 1187.540 1.120 1190.780 ;
  LAYER metal3 ;
  RECT 0.000 1187.540 1.120 1190.780 ;
  LAYER metal2 ;
  RECT 0.000 1187.540 1.120 1190.780 ;
  LAYER metal1 ;
  RECT 0.000 1187.540 1.120 1190.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1148.340 1.120 1151.580 ;
  LAYER metal4 ;
  RECT 0.000 1148.340 1.120 1151.580 ;
  LAYER metal3 ;
  RECT 0.000 1148.340 1.120 1151.580 ;
  LAYER metal2 ;
  RECT 0.000 1148.340 1.120 1151.580 ;
  LAYER metal1 ;
  RECT 0.000 1148.340 1.120 1151.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1140.500 1.120 1143.740 ;
  LAYER metal4 ;
  RECT 0.000 1140.500 1.120 1143.740 ;
  LAYER metal3 ;
  RECT 0.000 1140.500 1.120 1143.740 ;
  LAYER metal2 ;
  RECT 0.000 1140.500 1.120 1143.740 ;
  LAYER metal1 ;
  RECT 0.000 1140.500 1.120 1143.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1132.660 1.120 1135.900 ;
  LAYER metal4 ;
  RECT 0.000 1132.660 1.120 1135.900 ;
  LAYER metal3 ;
  RECT 0.000 1132.660 1.120 1135.900 ;
  LAYER metal2 ;
  RECT 0.000 1132.660 1.120 1135.900 ;
  LAYER metal1 ;
  RECT 0.000 1132.660 1.120 1135.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1124.820 1.120 1128.060 ;
  LAYER metal4 ;
  RECT 0.000 1124.820 1.120 1128.060 ;
  LAYER metal3 ;
  RECT 0.000 1124.820 1.120 1128.060 ;
  LAYER metal2 ;
  RECT 0.000 1124.820 1.120 1128.060 ;
  LAYER metal1 ;
  RECT 0.000 1124.820 1.120 1128.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1116.980 1.120 1120.220 ;
  LAYER metal4 ;
  RECT 0.000 1116.980 1.120 1120.220 ;
  LAYER metal3 ;
  RECT 0.000 1116.980 1.120 1120.220 ;
  LAYER metal2 ;
  RECT 0.000 1116.980 1.120 1120.220 ;
  LAYER metal1 ;
  RECT 0.000 1116.980 1.120 1120.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1109.140 1.120 1112.380 ;
  LAYER metal4 ;
  RECT 0.000 1109.140 1.120 1112.380 ;
  LAYER metal3 ;
  RECT 0.000 1109.140 1.120 1112.380 ;
  LAYER metal2 ;
  RECT 0.000 1109.140 1.120 1112.380 ;
  LAYER metal1 ;
  RECT 0.000 1109.140 1.120 1112.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1069.940 1.120 1073.180 ;
  LAYER metal4 ;
  RECT 0.000 1069.940 1.120 1073.180 ;
  LAYER metal3 ;
  RECT 0.000 1069.940 1.120 1073.180 ;
  LAYER metal2 ;
  RECT 0.000 1069.940 1.120 1073.180 ;
  LAYER metal1 ;
  RECT 0.000 1069.940 1.120 1073.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1062.100 1.120 1065.340 ;
  LAYER metal4 ;
  RECT 0.000 1062.100 1.120 1065.340 ;
  LAYER metal3 ;
  RECT 0.000 1062.100 1.120 1065.340 ;
  LAYER metal2 ;
  RECT 0.000 1062.100 1.120 1065.340 ;
  LAYER metal1 ;
  RECT 0.000 1062.100 1.120 1065.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1054.260 1.120 1057.500 ;
  LAYER metal4 ;
  RECT 0.000 1054.260 1.120 1057.500 ;
  LAYER metal3 ;
  RECT 0.000 1054.260 1.120 1057.500 ;
  LAYER metal2 ;
  RECT 0.000 1054.260 1.120 1057.500 ;
  LAYER metal1 ;
  RECT 0.000 1054.260 1.120 1057.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1046.420 1.120 1049.660 ;
  LAYER metal4 ;
  RECT 0.000 1046.420 1.120 1049.660 ;
  LAYER metal3 ;
  RECT 0.000 1046.420 1.120 1049.660 ;
  LAYER metal2 ;
  RECT 0.000 1046.420 1.120 1049.660 ;
  LAYER metal1 ;
  RECT 0.000 1046.420 1.120 1049.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1038.580 1.120 1041.820 ;
  LAYER metal4 ;
  RECT 0.000 1038.580 1.120 1041.820 ;
  LAYER metal3 ;
  RECT 0.000 1038.580 1.120 1041.820 ;
  LAYER metal2 ;
  RECT 0.000 1038.580 1.120 1041.820 ;
  LAYER metal1 ;
  RECT 0.000 1038.580 1.120 1041.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1030.740 1.120 1033.980 ;
  LAYER metal4 ;
  RECT 0.000 1030.740 1.120 1033.980 ;
  LAYER metal3 ;
  RECT 0.000 1030.740 1.120 1033.980 ;
  LAYER metal2 ;
  RECT 0.000 1030.740 1.120 1033.980 ;
  LAYER metal1 ;
  RECT 0.000 1030.740 1.120 1033.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 991.540 1.120 994.780 ;
  LAYER metal4 ;
  RECT 0.000 991.540 1.120 994.780 ;
  LAYER metal3 ;
  RECT 0.000 991.540 1.120 994.780 ;
  LAYER metal2 ;
  RECT 0.000 991.540 1.120 994.780 ;
  LAYER metal1 ;
  RECT 0.000 991.540 1.120 994.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 983.700 1.120 986.940 ;
  LAYER metal4 ;
  RECT 0.000 983.700 1.120 986.940 ;
  LAYER metal3 ;
  RECT 0.000 983.700 1.120 986.940 ;
  LAYER metal2 ;
  RECT 0.000 983.700 1.120 986.940 ;
  LAYER metal1 ;
  RECT 0.000 983.700 1.120 986.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 975.860 1.120 979.100 ;
  LAYER metal4 ;
  RECT 0.000 975.860 1.120 979.100 ;
  LAYER metal3 ;
  RECT 0.000 975.860 1.120 979.100 ;
  LAYER metal2 ;
  RECT 0.000 975.860 1.120 979.100 ;
  LAYER metal1 ;
  RECT 0.000 975.860 1.120 979.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 968.020 1.120 971.260 ;
  LAYER metal4 ;
  RECT 0.000 968.020 1.120 971.260 ;
  LAYER metal3 ;
  RECT 0.000 968.020 1.120 971.260 ;
  LAYER metal2 ;
  RECT 0.000 968.020 1.120 971.260 ;
  LAYER metal1 ;
  RECT 0.000 968.020 1.120 971.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 960.180 1.120 963.420 ;
  LAYER metal4 ;
  RECT 0.000 960.180 1.120 963.420 ;
  LAYER metal3 ;
  RECT 0.000 960.180 1.120 963.420 ;
  LAYER metal2 ;
  RECT 0.000 960.180 1.120 963.420 ;
  LAYER metal1 ;
  RECT 0.000 960.180 1.120 963.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 952.340 1.120 955.580 ;
  LAYER metal4 ;
  RECT 0.000 952.340 1.120 955.580 ;
  LAYER metal3 ;
  RECT 0.000 952.340 1.120 955.580 ;
  LAYER metal2 ;
  RECT 0.000 952.340 1.120 955.580 ;
  LAYER metal1 ;
  RECT 0.000 952.340 1.120 955.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 913.140 1.120 916.380 ;
  LAYER metal4 ;
  RECT 0.000 913.140 1.120 916.380 ;
  LAYER metal3 ;
  RECT 0.000 913.140 1.120 916.380 ;
  LAYER metal2 ;
  RECT 0.000 913.140 1.120 916.380 ;
  LAYER metal1 ;
  RECT 0.000 913.140 1.120 916.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 905.300 1.120 908.540 ;
  LAYER metal4 ;
  RECT 0.000 905.300 1.120 908.540 ;
  LAYER metal3 ;
  RECT 0.000 905.300 1.120 908.540 ;
  LAYER metal2 ;
  RECT 0.000 905.300 1.120 908.540 ;
  LAYER metal1 ;
  RECT 0.000 905.300 1.120 908.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 897.460 1.120 900.700 ;
  LAYER metal4 ;
  RECT 0.000 897.460 1.120 900.700 ;
  LAYER metal3 ;
  RECT 0.000 897.460 1.120 900.700 ;
  LAYER metal2 ;
  RECT 0.000 897.460 1.120 900.700 ;
  LAYER metal1 ;
  RECT 0.000 897.460 1.120 900.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 889.620 1.120 892.860 ;
  LAYER metal4 ;
  RECT 0.000 889.620 1.120 892.860 ;
  LAYER metal3 ;
  RECT 0.000 889.620 1.120 892.860 ;
  LAYER metal2 ;
  RECT 0.000 889.620 1.120 892.860 ;
  LAYER metal1 ;
  RECT 0.000 889.620 1.120 892.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 881.780 1.120 885.020 ;
  LAYER metal4 ;
  RECT 0.000 881.780 1.120 885.020 ;
  LAYER metal3 ;
  RECT 0.000 881.780 1.120 885.020 ;
  LAYER metal2 ;
  RECT 0.000 881.780 1.120 885.020 ;
  LAYER metal1 ;
  RECT 0.000 881.780 1.120 885.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 873.940 1.120 877.180 ;
  LAYER metal4 ;
  RECT 0.000 873.940 1.120 877.180 ;
  LAYER metal3 ;
  RECT 0.000 873.940 1.120 877.180 ;
  LAYER metal2 ;
  RECT 0.000 873.940 1.120 877.180 ;
  LAYER metal1 ;
  RECT 0.000 873.940 1.120 877.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 834.740 1.120 837.980 ;
  LAYER metal4 ;
  RECT 0.000 834.740 1.120 837.980 ;
  LAYER metal3 ;
  RECT 0.000 834.740 1.120 837.980 ;
  LAYER metal2 ;
  RECT 0.000 834.740 1.120 837.980 ;
  LAYER metal1 ;
  RECT 0.000 834.740 1.120 837.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 826.900 1.120 830.140 ;
  LAYER metal4 ;
  RECT 0.000 826.900 1.120 830.140 ;
  LAYER metal3 ;
  RECT 0.000 826.900 1.120 830.140 ;
  LAYER metal2 ;
  RECT 0.000 826.900 1.120 830.140 ;
  LAYER metal1 ;
  RECT 0.000 826.900 1.120 830.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 819.060 1.120 822.300 ;
  LAYER metal4 ;
  RECT 0.000 819.060 1.120 822.300 ;
  LAYER metal3 ;
  RECT 0.000 819.060 1.120 822.300 ;
  LAYER metal2 ;
  RECT 0.000 819.060 1.120 822.300 ;
  LAYER metal1 ;
  RECT 0.000 819.060 1.120 822.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 811.220 1.120 814.460 ;
  LAYER metal4 ;
  RECT 0.000 811.220 1.120 814.460 ;
  LAYER metal3 ;
  RECT 0.000 811.220 1.120 814.460 ;
  LAYER metal2 ;
  RECT 0.000 811.220 1.120 814.460 ;
  LAYER metal1 ;
  RECT 0.000 811.220 1.120 814.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 803.380 1.120 806.620 ;
  LAYER metal4 ;
  RECT 0.000 803.380 1.120 806.620 ;
  LAYER metal3 ;
  RECT 0.000 803.380 1.120 806.620 ;
  LAYER metal2 ;
  RECT 0.000 803.380 1.120 806.620 ;
  LAYER metal1 ;
  RECT 0.000 803.380 1.120 806.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 795.540 1.120 798.780 ;
  LAYER metal4 ;
  RECT 0.000 795.540 1.120 798.780 ;
  LAYER metal3 ;
  RECT 0.000 795.540 1.120 798.780 ;
  LAYER metal2 ;
  RECT 0.000 795.540 1.120 798.780 ;
  LAYER metal1 ;
  RECT 0.000 795.540 1.120 798.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 756.340 1.120 759.580 ;
  LAYER metal4 ;
  RECT 0.000 756.340 1.120 759.580 ;
  LAYER metal3 ;
  RECT 0.000 756.340 1.120 759.580 ;
  LAYER metal2 ;
  RECT 0.000 756.340 1.120 759.580 ;
  LAYER metal1 ;
  RECT 0.000 756.340 1.120 759.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 748.500 1.120 751.740 ;
  LAYER metal4 ;
  RECT 0.000 748.500 1.120 751.740 ;
  LAYER metal3 ;
  RECT 0.000 748.500 1.120 751.740 ;
  LAYER metal2 ;
  RECT 0.000 748.500 1.120 751.740 ;
  LAYER metal1 ;
  RECT 0.000 748.500 1.120 751.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 740.660 1.120 743.900 ;
  LAYER metal4 ;
  RECT 0.000 740.660 1.120 743.900 ;
  LAYER metal3 ;
  RECT 0.000 740.660 1.120 743.900 ;
  LAYER metal2 ;
  RECT 0.000 740.660 1.120 743.900 ;
  LAYER metal1 ;
  RECT 0.000 740.660 1.120 743.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 732.820 1.120 736.060 ;
  LAYER metal4 ;
  RECT 0.000 732.820 1.120 736.060 ;
  LAYER metal3 ;
  RECT 0.000 732.820 1.120 736.060 ;
  LAYER metal2 ;
  RECT 0.000 732.820 1.120 736.060 ;
  LAYER metal1 ;
  RECT 0.000 732.820 1.120 736.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 724.980 1.120 728.220 ;
  LAYER metal4 ;
  RECT 0.000 724.980 1.120 728.220 ;
  LAYER metal3 ;
  RECT 0.000 724.980 1.120 728.220 ;
  LAYER metal2 ;
  RECT 0.000 724.980 1.120 728.220 ;
  LAYER metal1 ;
  RECT 0.000 724.980 1.120 728.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 717.140 1.120 720.380 ;
  LAYER metal4 ;
  RECT 0.000 717.140 1.120 720.380 ;
  LAYER metal3 ;
  RECT 0.000 717.140 1.120 720.380 ;
  LAYER metal2 ;
  RECT 0.000 717.140 1.120 720.380 ;
  LAYER metal1 ;
  RECT 0.000 717.140 1.120 720.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 677.940 1.120 681.180 ;
  LAYER metal4 ;
  RECT 0.000 677.940 1.120 681.180 ;
  LAYER metal3 ;
  RECT 0.000 677.940 1.120 681.180 ;
  LAYER metal2 ;
  RECT 0.000 677.940 1.120 681.180 ;
  LAYER metal1 ;
  RECT 0.000 677.940 1.120 681.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 670.100 1.120 673.340 ;
  LAYER metal4 ;
  RECT 0.000 670.100 1.120 673.340 ;
  LAYER metal3 ;
  RECT 0.000 670.100 1.120 673.340 ;
  LAYER metal2 ;
  RECT 0.000 670.100 1.120 673.340 ;
  LAYER metal1 ;
  RECT 0.000 670.100 1.120 673.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 662.260 1.120 665.500 ;
  LAYER metal4 ;
  RECT 0.000 662.260 1.120 665.500 ;
  LAYER metal3 ;
  RECT 0.000 662.260 1.120 665.500 ;
  LAYER metal2 ;
  RECT 0.000 662.260 1.120 665.500 ;
  LAYER metal1 ;
  RECT 0.000 662.260 1.120 665.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 654.420 1.120 657.660 ;
  LAYER metal4 ;
  RECT 0.000 654.420 1.120 657.660 ;
  LAYER metal3 ;
  RECT 0.000 654.420 1.120 657.660 ;
  LAYER metal2 ;
  RECT 0.000 654.420 1.120 657.660 ;
  LAYER metal1 ;
  RECT 0.000 654.420 1.120 657.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 646.580 1.120 649.820 ;
  LAYER metal4 ;
  RECT 0.000 646.580 1.120 649.820 ;
  LAYER metal3 ;
  RECT 0.000 646.580 1.120 649.820 ;
  LAYER metal2 ;
  RECT 0.000 646.580 1.120 649.820 ;
  LAYER metal1 ;
  RECT 0.000 646.580 1.120 649.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 638.740 1.120 641.980 ;
  LAYER metal4 ;
  RECT 0.000 638.740 1.120 641.980 ;
  LAYER metal3 ;
  RECT 0.000 638.740 1.120 641.980 ;
  LAYER metal2 ;
  RECT 0.000 638.740 1.120 641.980 ;
  LAYER metal1 ;
  RECT 0.000 638.740 1.120 641.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 599.540 1.120 602.780 ;
  LAYER metal4 ;
  RECT 0.000 599.540 1.120 602.780 ;
  LAYER metal3 ;
  RECT 0.000 599.540 1.120 602.780 ;
  LAYER metal2 ;
  RECT 0.000 599.540 1.120 602.780 ;
  LAYER metal1 ;
  RECT 0.000 599.540 1.120 602.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 591.700 1.120 594.940 ;
  LAYER metal4 ;
  RECT 0.000 591.700 1.120 594.940 ;
  LAYER metal3 ;
  RECT 0.000 591.700 1.120 594.940 ;
  LAYER metal2 ;
  RECT 0.000 591.700 1.120 594.940 ;
  LAYER metal1 ;
  RECT 0.000 591.700 1.120 594.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 583.860 1.120 587.100 ;
  LAYER metal4 ;
  RECT 0.000 583.860 1.120 587.100 ;
  LAYER metal3 ;
  RECT 0.000 583.860 1.120 587.100 ;
  LAYER metal2 ;
  RECT 0.000 583.860 1.120 587.100 ;
  LAYER metal1 ;
  RECT 0.000 583.860 1.120 587.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 576.020 1.120 579.260 ;
  LAYER metal4 ;
  RECT 0.000 576.020 1.120 579.260 ;
  LAYER metal3 ;
  RECT 0.000 576.020 1.120 579.260 ;
  LAYER metal2 ;
  RECT 0.000 576.020 1.120 579.260 ;
  LAYER metal1 ;
  RECT 0.000 576.020 1.120 579.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 568.180 1.120 571.420 ;
  LAYER metal4 ;
  RECT 0.000 568.180 1.120 571.420 ;
  LAYER metal3 ;
  RECT 0.000 568.180 1.120 571.420 ;
  LAYER metal2 ;
  RECT 0.000 568.180 1.120 571.420 ;
  LAYER metal1 ;
  RECT 0.000 568.180 1.120 571.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 560.340 1.120 563.580 ;
  LAYER metal4 ;
  RECT 0.000 560.340 1.120 563.580 ;
  LAYER metal3 ;
  RECT 0.000 560.340 1.120 563.580 ;
  LAYER metal2 ;
  RECT 0.000 560.340 1.120 563.580 ;
  LAYER metal1 ;
  RECT 0.000 560.340 1.120 563.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 521.140 1.120 524.380 ;
  LAYER metal4 ;
  RECT 0.000 521.140 1.120 524.380 ;
  LAYER metal3 ;
  RECT 0.000 521.140 1.120 524.380 ;
  LAYER metal2 ;
  RECT 0.000 521.140 1.120 524.380 ;
  LAYER metal1 ;
  RECT 0.000 521.140 1.120 524.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 513.300 1.120 516.540 ;
  LAYER metal4 ;
  RECT 0.000 513.300 1.120 516.540 ;
  LAYER metal3 ;
  RECT 0.000 513.300 1.120 516.540 ;
  LAYER metal2 ;
  RECT 0.000 513.300 1.120 516.540 ;
  LAYER metal1 ;
  RECT 0.000 513.300 1.120 516.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 505.460 1.120 508.700 ;
  LAYER metal4 ;
  RECT 0.000 505.460 1.120 508.700 ;
  LAYER metal3 ;
  RECT 0.000 505.460 1.120 508.700 ;
  LAYER metal2 ;
  RECT 0.000 505.460 1.120 508.700 ;
  LAYER metal1 ;
  RECT 0.000 505.460 1.120 508.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 497.620 1.120 500.860 ;
  LAYER metal4 ;
  RECT 0.000 497.620 1.120 500.860 ;
  LAYER metal3 ;
  RECT 0.000 497.620 1.120 500.860 ;
  LAYER metal2 ;
  RECT 0.000 497.620 1.120 500.860 ;
  LAYER metal1 ;
  RECT 0.000 497.620 1.120 500.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 489.780 1.120 493.020 ;
  LAYER metal4 ;
  RECT 0.000 489.780 1.120 493.020 ;
  LAYER metal3 ;
  RECT 0.000 489.780 1.120 493.020 ;
  LAYER metal2 ;
  RECT 0.000 489.780 1.120 493.020 ;
  LAYER metal1 ;
  RECT 0.000 489.780 1.120 493.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 481.940 1.120 485.180 ;
  LAYER metal4 ;
  RECT 0.000 481.940 1.120 485.180 ;
  LAYER metal3 ;
  RECT 0.000 481.940 1.120 485.180 ;
  LAYER metal2 ;
  RECT 0.000 481.940 1.120 485.180 ;
  LAYER metal1 ;
  RECT 0.000 481.940 1.120 485.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 442.740 1.120 445.980 ;
  LAYER metal4 ;
  RECT 0.000 442.740 1.120 445.980 ;
  LAYER metal3 ;
  RECT 0.000 442.740 1.120 445.980 ;
  LAYER metal2 ;
  RECT 0.000 442.740 1.120 445.980 ;
  LAYER metal1 ;
  RECT 0.000 442.740 1.120 445.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 434.900 1.120 438.140 ;
  LAYER metal4 ;
  RECT 0.000 434.900 1.120 438.140 ;
  LAYER metal3 ;
  RECT 0.000 434.900 1.120 438.140 ;
  LAYER metal2 ;
  RECT 0.000 434.900 1.120 438.140 ;
  LAYER metal1 ;
  RECT 0.000 434.900 1.120 438.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 427.060 1.120 430.300 ;
  LAYER metal4 ;
  RECT 0.000 427.060 1.120 430.300 ;
  LAYER metal3 ;
  RECT 0.000 427.060 1.120 430.300 ;
  LAYER metal2 ;
  RECT 0.000 427.060 1.120 430.300 ;
  LAYER metal1 ;
  RECT 0.000 427.060 1.120 430.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 419.220 1.120 422.460 ;
  LAYER metal4 ;
  RECT 0.000 419.220 1.120 422.460 ;
  LAYER metal3 ;
  RECT 0.000 419.220 1.120 422.460 ;
  LAYER metal2 ;
  RECT 0.000 419.220 1.120 422.460 ;
  LAYER metal1 ;
  RECT 0.000 419.220 1.120 422.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 411.380 1.120 414.620 ;
  LAYER metal4 ;
  RECT 0.000 411.380 1.120 414.620 ;
  LAYER metal3 ;
  RECT 0.000 411.380 1.120 414.620 ;
  LAYER metal2 ;
  RECT 0.000 411.380 1.120 414.620 ;
  LAYER metal1 ;
  RECT 0.000 411.380 1.120 414.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 403.540 1.120 406.780 ;
  LAYER metal4 ;
  RECT 0.000 403.540 1.120 406.780 ;
  LAYER metal3 ;
  RECT 0.000 403.540 1.120 406.780 ;
  LAYER metal2 ;
  RECT 0.000 403.540 1.120 406.780 ;
  LAYER metal1 ;
  RECT 0.000 403.540 1.120 406.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 364.340 1.120 367.580 ;
  LAYER metal4 ;
  RECT 0.000 364.340 1.120 367.580 ;
  LAYER metal3 ;
  RECT 0.000 364.340 1.120 367.580 ;
  LAYER metal2 ;
  RECT 0.000 364.340 1.120 367.580 ;
  LAYER metal1 ;
  RECT 0.000 364.340 1.120 367.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 356.500 1.120 359.740 ;
  LAYER metal4 ;
  RECT 0.000 356.500 1.120 359.740 ;
  LAYER metal3 ;
  RECT 0.000 356.500 1.120 359.740 ;
  LAYER metal2 ;
  RECT 0.000 356.500 1.120 359.740 ;
  LAYER metal1 ;
  RECT 0.000 356.500 1.120 359.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 348.660 1.120 351.900 ;
  LAYER metal4 ;
  RECT 0.000 348.660 1.120 351.900 ;
  LAYER metal3 ;
  RECT 0.000 348.660 1.120 351.900 ;
  LAYER metal2 ;
  RECT 0.000 348.660 1.120 351.900 ;
  LAYER metal1 ;
  RECT 0.000 348.660 1.120 351.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 340.820 1.120 344.060 ;
  LAYER metal4 ;
  RECT 0.000 340.820 1.120 344.060 ;
  LAYER metal3 ;
  RECT 0.000 340.820 1.120 344.060 ;
  LAYER metal2 ;
  RECT 0.000 340.820 1.120 344.060 ;
  LAYER metal1 ;
  RECT 0.000 340.820 1.120 344.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 332.980 1.120 336.220 ;
  LAYER metal4 ;
  RECT 0.000 332.980 1.120 336.220 ;
  LAYER metal3 ;
  RECT 0.000 332.980 1.120 336.220 ;
  LAYER metal2 ;
  RECT 0.000 332.980 1.120 336.220 ;
  LAYER metal1 ;
  RECT 0.000 332.980 1.120 336.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 325.140 1.120 328.380 ;
  LAYER metal4 ;
  RECT 0.000 325.140 1.120 328.380 ;
  LAYER metal3 ;
  RECT 0.000 325.140 1.120 328.380 ;
  LAYER metal2 ;
  RECT 0.000 325.140 1.120 328.380 ;
  LAYER metal1 ;
  RECT 0.000 325.140 1.120 328.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 285.940 1.120 289.180 ;
  LAYER metal4 ;
  RECT 0.000 285.940 1.120 289.180 ;
  LAYER metal3 ;
  RECT 0.000 285.940 1.120 289.180 ;
  LAYER metal2 ;
  RECT 0.000 285.940 1.120 289.180 ;
  LAYER metal1 ;
  RECT 0.000 285.940 1.120 289.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 278.100 1.120 281.340 ;
  LAYER metal4 ;
  RECT 0.000 278.100 1.120 281.340 ;
  LAYER metal3 ;
  RECT 0.000 278.100 1.120 281.340 ;
  LAYER metal2 ;
  RECT 0.000 278.100 1.120 281.340 ;
  LAYER metal1 ;
  RECT 0.000 278.100 1.120 281.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 270.260 1.120 273.500 ;
  LAYER metal4 ;
  RECT 0.000 270.260 1.120 273.500 ;
  LAYER metal3 ;
  RECT 0.000 270.260 1.120 273.500 ;
  LAYER metal2 ;
  RECT 0.000 270.260 1.120 273.500 ;
  LAYER metal1 ;
  RECT 0.000 270.260 1.120 273.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 262.420 1.120 265.660 ;
  LAYER metal4 ;
  RECT 0.000 262.420 1.120 265.660 ;
  LAYER metal3 ;
  RECT 0.000 262.420 1.120 265.660 ;
  LAYER metal2 ;
  RECT 0.000 262.420 1.120 265.660 ;
  LAYER metal1 ;
  RECT 0.000 262.420 1.120 265.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 254.580 1.120 257.820 ;
  LAYER metal4 ;
  RECT 0.000 254.580 1.120 257.820 ;
  LAYER metal3 ;
  RECT 0.000 254.580 1.120 257.820 ;
  LAYER metal2 ;
  RECT 0.000 254.580 1.120 257.820 ;
  LAYER metal1 ;
  RECT 0.000 254.580 1.120 257.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 246.740 1.120 249.980 ;
  LAYER metal4 ;
  RECT 0.000 246.740 1.120 249.980 ;
  LAYER metal3 ;
  RECT 0.000 246.740 1.120 249.980 ;
  LAYER metal2 ;
  RECT 0.000 246.740 1.120 249.980 ;
  LAYER metal1 ;
  RECT 0.000 246.740 1.120 249.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 207.540 1.120 210.780 ;
  LAYER metal4 ;
  RECT 0.000 207.540 1.120 210.780 ;
  LAYER metal3 ;
  RECT 0.000 207.540 1.120 210.780 ;
  LAYER metal2 ;
  RECT 0.000 207.540 1.120 210.780 ;
  LAYER metal1 ;
  RECT 0.000 207.540 1.120 210.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER metal4 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER metal3 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER metal2 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER metal1 ;
  RECT 0.000 199.700 1.120 202.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER metal4 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER metal3 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER metal2 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER metal1 ;
  RECT 0.000 191.860 1.120 195.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER metal4 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER metal3 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER metal2 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER metal1 ;
  RECT 0.000 184.020 1.120 187.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER metal4 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER metal3 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER metal2 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER metal1 ;
  RECT 0.000 176.180 1.120 179.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER metal4 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER metal3 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER metal2 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER metal1 ;
  RECT 0.000 168.340 1.120 171.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER metal4 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER metal3 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER metal2 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER metal1 ;
  RECT 0.000 129.140 1.120 132.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER metal4 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER metal3 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER metal2 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER metal1 ;
  RECT 0.000 121.300 1.120 124.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER metal4 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER metal3 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER metal2 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER metal1 ;
  RECT 0.000 113.460 1.120 116.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER metal4 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER metal3 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER metal2 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER metal1 ;
  RECT 0.000 105.620 1.120 108.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER metal4 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER metal3 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER metal2 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER metal1 ;
  RECT 0.000 97.780 1.120 101.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER metal4 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER metal3 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER metal2 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER metal1 ;
  RECT 0.000 89.940 1.120 93.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER metal4 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER metal3 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER metal2 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER metal1 ;
  RECT 0.000 50.740 1.120 53.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER metal4 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER metal3 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER metal2 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER metal1 ;
  RECT 0.000 42.900 1.120 46.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER metal4 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER metal3 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER metal2 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER metal1 ;
  RECT 0.000 35.060 1.120 38.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER metal4 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER metal3 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER metal2 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER metal1 ;
  RECT 0.000 27.220 1.120 30.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER metal4 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER metal3 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER metal2 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER metal1 ;
  RECT 0.000 19.380 1.120 22.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER metal4 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER metal3 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER metal2 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER metal1 ;
  RECT 0.000 11.540 1.120 14.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3592.060 1710.800 3595.600 1711.920 ;
  LAYER metal4 ;
  RECT 3592.060 1710.800 3595.600 1711.920 ;
  LAYER metal3 ;
  RECT 3592.060 1710.800 3595.600 1711.920 ;
  LAYER metal2 ;
  RECT 3592.060 1710.800 3595.600 1711.920 ;
  LAYER metal1 ;
  RECT 3592.060 1710.800 3595.600 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3583.380 1710.800 3586.920 1711.920 ;
  LAYER metal4 ;
  RECT 3583.380 1710.800 3586.920 1711.920 ;
  LAYER metal3 ;
  RECT 3583.380 1710.800 3586.920 1711.920 ;
  LAYER metal2 ;
  RECT 3583.380 1710.800 3586.920 1711.920 ;
  LAYER metal1 ;
  RECT 3583.380 1710.800 3586.920 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3574.700 1710.800 3578.240 1711.920 ;
  LAYER metal4 ;
  RECT 3574.700 1710.800 3578.240 1711.920 ;
  LAYER metal3 ;
  RECT 3574.700 1710.800 3578.240 1711.920 ;
  LAYER metal2 ;
  RECT 3574.700 1710.800 3578.240 1711.920 ;
  LAYER metal1 ;
  RECT 3574.700 1710.800 3578.240 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3566.020 1710.800 3569.560 1711.920 ;
  LAYER metal4 ;
  RECT 3566.020 1710.800 3569.560 1711.920 ;
  LAYER metal3 ;
  RECT 3566.020 1710.800 3569.560 1711.920 ;
  LAYER metal2 ;
  RECT 3566.020 1710.800 3569.560 1711.920 ;
  LAYER metal1 ;
  RECT 3566.020 1710.800 3569.560 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3557.340 1710.800 3560.880 1711.920 ;
  LAYER metal4 ;
  RECT 3557.340 1710.800 3560.880 1711.920 ;
  LAYER metal3 ;
  RECT 3557.340 1710.800 3560.880 1711.920 ;
  LAYER metal2 ;
  RECT 3557.340 1710.800 3560.880 1711.920 ;
  LAYER metal1 ;
  RECT 3557.340 1710.800 3560.880 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3548.660 1710.800 3552.200 1711.920 ;
  LAYER metal4 ;
  RECT 3548.660 1710.800 3552.200 1711.920 ;
  LAYER metal3 ;
  RECT 3548.660 1710.800 3552.200 1711.920 ;
  LAYER metal2 ;
  RECT 3548.660 1710.800 3552.200 1711.920 ;
  LAYER metal1 ;
  RECT 3548.660 1710.800 3552.200 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3505.260 1710.800 3508.800 1711.920 ;
  LAYER metal4 ;
  RECT 3505.260 1710.800 3508.800 1711.920 ;
  LAYER metal3 ;
  RECT 3505.260 1710.800 3508.800 1711.920 ;
  LAYER metal2 ;
  RECT 3505.260 1710.800 3508.800 1711.920 ;
  LAYER metal1 ;
  RECT 3505.260 1710.800 3508.800 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3496.580 1710.800 3500.120 1711.920 ;
  LAYER metal4 ;
  RECT 3496.580 1710.800 3500.120 1711.920 ;
  LAYER metal3 ;
  RECT 3496.580 1710.800 3500.120 1711.920 ;
  LAYER metal2 ;
  RECT 3496.580 1710.800 3500.120 1711.920 ;
  LAYER metal1 ;
  RECT 3496.580 1710.800 3500.120 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3487.900 1710.800 3491.440 1711.920 ;
  LAYER metal4 ;
  RECT 3487.900 1710.800 3491.440 1711.920 ;
  LAYER metal3 ;
  RECT 3487.900 1710.800 3491.440 1711.920 ;
  LAYER metal2 ;
  RECT 3487.900 1710.800 3491.440 1711.920 ;
  LAYER metal1 ;
  RECT 3487.900 1710.800 3491.440 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3479.220 1710.800 3482.760 1711.920 ;
  LAYER metal4 ;
  RECT 3479.220 1710.800 3482.760 1711.920 ;
  LAYER metal3 ;
  RECT 3479.220 1710.800 3482.760 1711.920 ;
  LAYER metal2 ;
  RECT 3479.220 1710.800 3482.760 1711.920 ;
  LAYER metal1 ;
  RECT 3479.220 1710.800 3482.760 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3470.540 1710.800 3474.080 1711.920 ;
  LAYER metal4 ;
  RECT 3470.540 1710.800 3474.080 1711.920 ;
  LAYER metal3 ;
  RECT 3470.540 1710.800 3474.080 1711.920 ;
  LAYER metal2 ;
  RECT 3470.540 1710.800 3474.080 1711.920 ;
  LAYER metal1 ;
  RECT 3470.540 1710.800 3474.080 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3461.860 1710.800 3465.400 1711.920 ;
  LAYER metal4 ;
  RECT 3461.860 1710.800 3465.400 1711.920 ;
  LAYER metal3 ;
  RECT 3461.860 1710.800 3465.400 1711.920 ;
  LAYER metal2 ;
  RECT 3461.860 1710.800 3465.400 1711.920 ;
  LAYER metal1 ;
  RECT 3461.860 1710.800 3465.400 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3418.460 1710.800 3422.000 1711.920 ;
  LAYER metal4 ;
  RECT 3418.460 1710.800 3422.000 1711.920 ;
  LAYER metal3 ;
  RECT 3418.460 1710.800 3422.000 1711.920 ;
  LAYER metal2 ;
  RECT 3418.460 1710.800 3422.000 1711.920 ;
  LAYER metal1 ;
  RECT 3418.460 1710.800 3422.000 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3409.780 1710.800 3413.320 1711.920 ;
  LAYER metal4 ;
  RECT 3409.780 1710.800 3413.320 1711.920 ;
  LAYER metal3 ;
  RECT 3409.780 1710.800 3413.320 1711.920 ;
  LAYER metal2 ;
  RECT 3409.780 1710.800 3413.320 1711.920 ;
  LAYER metal1 ;
  RECT 3409.780 1710.800 3413.320 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3401.100 1710.800 3404.640 1711.920 ;
  LAYER metal4 ;
  RECT 3401.100 1710.800 3404.640 1711.920 ;
  LAYER metal3 ;
  RECT 3401.100 1710.800 3404.640 1711.920 ;
  LAYER metal2 ;
  RECT 3401.100 1710.800 3404.640 1711.920 ;
  LAYER metal1 ;
  RECT 3401.100 1710.800 3404.640 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3392.420 1710.800 3395.960 1711.920 ;
  LAYER metal4 ;
  RECT 3392.420 1710.800 3395.960 1711.920 ;
  LAYER metal3 ;
  RECT 3392.420 1710.800 3395.960 1711.920 ;
  LAYER metal2 ;
  RECT 3392.420 1710.800 3395.960 1711.920 ;
  LAYER metal1 ;
  RECT 3392.420 1710.800 3395.960 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3383.740 1710.800 3387.280 1711.920 ;
  LAYER metal4 ;
  RECT 3383.740 1710.800 3387.280 1711.920 ;
  LAYER metal3 ;
  RECT 3383.740 1710.800 3387.280 1711.920 ;
  LAYER metal2 ;
  RECT 3383.740 1710.800 3387.280 1711.920 ;
  LAYER metal1 ;
  RECT 3383.740 1710.800 3387.280 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3375.060 1710.800 3378.600 1711.920 ;
  LAYER metal4 ;
  RECT 3375.060 1710.800 3378.600 1711.920 ;
  LAYER metal3 ;
  RECT 3375.060 1710.800 3378.600 1711.920 ;
  LAYER metal2 ;
  RECT 3375.060 1710.800 3378.600 1711.920 ;
  LAYER metal1 ;
  RECT 3375.060 1710.800 3378.600 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3331.660 1710.800 3335.200 1711.920 ;
  LAYER metal4 ;
  RECT 3331.660 1710.800 3335.200 1711.920 ;
  LAYER metal3 ;
  RECT 3331.660 1710.800 3335.200 1711.920 ;
  LAYER metal2 ;
  RECT 3331.660 1710.800 3335.200 1711.920 ;
  LAYER metal1 ;
  RECT 3331.660 1710.800 3335.200 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3322.980 1710.800 3326.520 1711.920 ;
  LAYER metal4 ;
  RECT 3322.980 1710.800 3326.520 1711.920 ;
  LAYER metal3 ;
  RECT 3322.980 1710.800 3326.520 1711.920 ;
  LAYER metal2 ;
  RECT 3322.980 1710.800 3326.520 1711.920 ;
  LAYER metal1 ;
  RECT 3322.980 1710.800 3326.520 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3314.300 1710.800 3317.840 1711.920 ;
  LAYER metal4 ;
  RECT 3314.300 1710.800 3317.840 1711.920 ;
  LAYER metal3 ;
  RECT 3314.300 1710.800 3317.840 1711.920 ;
  LAYER metal2 ;
  RECT 3314.300 1710.800 3317.840 1711.920 ;
  LAYER metal1 ;
  RECT 3314.300 1710.800 3317.840 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3305.620 1710.800 3309.160 1711.920 ;
  LAYER metal4 ;
  RECT 3305.620 1710.800 3309.160 1711.920 ;
  LAYER metal3 ;
  RECT 3305.620 1710.800 3309.160 1711.920 ;
  LAYER metal2 ;
  RECT 3305.620 1710.800 3309.160 1711.920 ;
  LAYER metal1 ;
  RECT 3305.620 1710.800 3309.160 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3296.940 1710.800 3300.480 1711.920 ;
  LAYER metal4 ;
  RECT 3296.940 1710.800 3300.480 1711.920 ;
  LAYER metal3 ;
  RECT 3296.940 1710.800 3300.480 1711.920 ;
  LAYER metal2 ;
  RECT 3296.940 1710.800 3300.480 1711.920 ;
  LAYER metal1 ;
  RECT 3296.940 1710.800 3300.480 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3288.260 1710.800 3291.800 1711.920 ;
  LAYER metal4 ;
  RECT 3288.260 1710.800 3291.800 1711.920 ;
  LAYER metal3 ;
  RECT 3288.260 1710.800 3291.800 1711.920 ;
  LAYER metal2 ;
  RECT 3288.260 1710.800 3291.800 1711.920 ;
  LAYER metal1 ;
  RECT 3288.260 1710.800 3291.800 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3244.860 1710.800 3248.400 1711.920 ;
  LAYER metal4 ;
  RECT 3244.860 1710.800 3248.400 1711.920 ;
  LAYER metal3 ;
  RECT 3244.860 1710.800 3248.400 1711.920 ;
  LAYER metal2 ;
  RECT 3244.860 1710.800 3248.400 1711.920 ;
  LAYER metal1 ;
  RECT 3244.860 1710.800 3248.400 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3236.180 1710.800 3239.720 1711.920 ;
  LAYER metal4 ;
  RECT 3236.180 1710.800 3239.720 1711.920 ;
  LAYER metal3 ;
  RECT 3236.180 1710.800 3239.720 1711.920 ;
  LAYER metal2 ;
  RECT 3236.180 1710.800 3239.720 1711.920 ;
  LAYER metal1 ;
  RECT 3236.180 1710.800 3239.720 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3227.500 1710.800 3231.040 1711.920 ;
  LAYER metal4 ;
  RECT 3227.500 1710.800 3231.040 1711.920 ;
  LAYER metal3 ;
  RECT 3227.500 1710.800 3231.040 1711.920 ;
  LAYER metal2 ;
  RECT 3227.500 1710.800 3231.040 1711.920 ;
  LAYER metal1 ;
  RECT 3227.500 1710.800 3231.040 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3218.820 1710.800 3222.360 1711.920 ;
  LAYER metal4 ;
  RECT 3218.820 1710.800 3222.360 1711.920 ;
  LAYER metal3 ;
  RECT 3218.820 1710.800 3222.360 1711.920 ;
  LAYER metal2 ;
  RECT 3218.820 1710.800 3222.360 1711.920 ;
  LAYER metal1 ;
  RECT 3218.820 1710.800 3222.360 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3205.800 1710.800 3209.340 1711.920 ;
  LAYER metal4 ;
  RECT 3205.800 1710.800 3209.340 1711.920 ;
  LAYER metal3 ;
  RECT 3205.800 1710.800 3209.340 1711.920 ;
  LAYER metal2 ;
  RECT 3205.800 1710.800 3209.340 1711.920 ;
  LAYER metal1 ;
  RECT 3205.800 1710.800 3209.340 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3192.160 1710.800 3195.700 1711.920 ;
  LAYER metal4 ;
  RECT 3192.160 1710.800 3195.700 1711.920 ;
  LAYER metal3 ;
  RECT 3192.160 1710.800 3195.700 1711.920 ;
  LAYER metal2 ;
  RECT 3192.160 1710.800 3195.700 1711.920 ;
  LAYER metal1 ;
  RECT 3192.160 1710.800 3195.700 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3138.220 1710.800 3141.760 1711.920 ;
  LAYER metal4 ;
  RECT 3138.220 1710.800 3141.760 1711.920 ;
  LAYER metal3 ;
  RECT 3138.220 1710.800 3141.760 1711.920 ;
  LAYER metal2 ;
  RECT 3138.220 1710.800 3141.760 1711.920 ;
  LAYER metal1 ;
  RECT 3138.220 1710.800 3141.760 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3129.540 1710.800 3133.080 1711.920 ;
  LAYER metal4 ;
  RECT 3129.540 1710.800 3133.080 1711.920 ;
  LAYER metal3 ;
  RECT 3129.540 1710.800 3133.080 1711.920 ;
  LAYER metal2 ;
  RECT 3129.540 1710.800 3133.080 1711.920 ;
  LAYER metal1 ;
  RECT 3129.540 1710.800 3133.080 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3120.860 1710.800 3124.400 1711.920 ;
  LAYER metal4 ;
  RECT 3120.860 1710.800 3124.400 1711.920 ;
  LAYER metal3 ;
  RECT 3120.860 1710.800 3124.400 1711.920 ;
  LAYER metal2 ;
  RECT 3120.860 1710.800 3124.400 1711.920 ;
  LAYER metal1 ;
  RECT 3120.860 1710.800 3124.400 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3112.180 1710.800 3115.720 1711.920 ;
  LAYER metal4 ;
  RECT 3112.180 1710.800 3115.720 1711.920 ;
  LAYER metal3 ;
  RECT 3112.180 1710.800 3115.720 1711.920 ;
  LAYER metal2 ;
  RECT 3112.180 1710.800 3115.720 1711.920 ;
  LAYER metal1 ;
  RECT 3112.180 1710.800 3115.720 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3103.500 1710.800 3107.040 1711.920 ;
  LAYER metal4 ;
  RECT 3103.500 1710.800 3107.040 1711.920 ;
  LAYER metal3 ;
  RECT 3103.500 1710.800 3107.040 1711.920 ;
  LAYER metal2 ;
  RECT 3103.500 1710.800 3107.040 1711.920 ;
  LAYER metal1 ;
  RECT 3103.500 1710.800 3107.040 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3094.820 1710.800 3098.360 1711.920 ;
  LAYER metal4 ;
  RECT 3094.820 1710.800 3098.360 1711.920 ;
  LAYER metal3 ;
  RECT 3094.820 1710.800 3098.360 1711.920 ;
  LAYER metal2 ;
  RECT 3094.820 1710.800 3098.360 1711.920 ;
  LAYER metal1 ;
  RECT 3094.820 1710.800 3098.360 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3051.420 1710.800 3054.960 1711.920 ;
  LAYER metal4 ;
  RECT 3051.420 1710.800 3054.960 1711.920 ;
  LAYER metal3 ;
  RECT 3051.420 1710.800 3054.960 1711.920 ;
  LAYER metal2 ;
  RECT 3051.420 1710.800 3054.960 1711.920 ;
  LAYER metal1 ;
  RECT 3051.420 1710.800 3054.960 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3042.740 1710.800 3046.280 1711.920 ;
  LAYER metal4 ;
  RECT 3042.740 1710.800 3046.280 1711.920 ;
  LAYER metal3 ;
  RECT 3042.740 1710.800 3046.280 1711.920 ;
  LAYER metal2 ;
  RECT 3042.740 1710.800 3046.280 1711.920 ;
  LAYER metal1 ;
  RECT 3042.740 1710.800 3046.280 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3034.060 1710.800 3037.600 1711.920 ;
  LAYER metal4 ;
  RECT 3034.060 1710.800 3037.600 1711.920 ;
  LAYER metal3 ;
  RECT 3034.060 1710.800 3037.600 1711.920 ;
  LAYER metal2 ;
  RECT 3034.060 1710.800 3037.600 1711.920 ;
  LAYER metal1 ;
  RECT 3034.060 1710.800 3037.600 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3025.380 1710.800 3028.920 1711.920 ;
  LAYER metal4 ;
  RECT 3025.380 1710.800 3028.920 1711.920 ;
  LAYER metal3 ;
  RECT 3025.380 1710.800 3028.920 1711.920 ;
  LAYER metal2 ;
  RECT 3025.380 1710.800 3028.920 1711.920 ;
  LAYER metal1 ;
  RECT 3025.380 1710.800 3028.920 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3016.700 1710.800 3020.240 1711.920 ;
  LAYER metal4 ;
  RECT 3016.700 1710.800 3020.240 1711.920 ;
  LAYER metal3 ;
  RECT 3016.700 1710.800 3020.240 1711.920 ;
  LAYER metal2 ;
  RECT 3016.700 1710.800 3020.240 1711.920 ;
  LAYER metal1 ;
  RECT 3016.700 1710.800 3020.240 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3008.020 1710.800 3011.560 1711.920 ;
  LAYER metal4 ;
  RECT 3008.020 1710.800 3011.560 1711.920 ;
  LAYER metal3 ;
  RECT 3008.020 1710.800 3011.560 1711.920 ;
  LAYER metal2 ;
  RECT 3008.020 1710.800 3011.560 1711.920 ;
  LAYER metal1 ;
  RECT 3008.020 1710.800 3011.560 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2964.620 1710.800 2968.160 1711.920 ;
  LAYER metal4 ;
  RECT 2964.620 1710.800 2968.160 1711.920 ;
  LAYER metal3 ;
  RECT 2964.620 1710.800 2968.160 1711.920 ;
  LAYER metal2 ;
  RECT 2964.620 1710.800 2968.160 1711.920 ;
  LAYER metal1 ;
  RECT 2964.620 1710.800 2968.160 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2955.940 1710.800 2959.480 1711.920 ;
  LAYER metal4 ;
  RECT 2955.940 1710.800 2959.480 1711.920 ;
  LAYER metal3 ;
  RECT 2955.940 1710.800 2959.480 1711.920 ;
  LAYER metal2 ;
  RECT 2955.940 1710.800 2959.480 1711.920 ;
  LAYER metal1 ;
  RECT 2955.940 1710.800 2959.480 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2947.260 1710.800 2950.800 1711.920 ;
  LAYER metal4 ;
  RECT 2947.260 1710.800 2950.800 1711.920 ;
  LAYER metal3 ;
  RECT 2947.260 1710.800 2950.800 1711.920 ;
  LAYER metal2 ;
  RECT 2947.260 1710.800 2950.800 1711.920 ;
  LAYER metal1 ;
  RECT 2947.260 1710.800 2950.800 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2938.580 1710.800 2942.120 1711.920 ;
  LAYER metal4 ;
  RECT 2938.580 1710.800 2942.120 1711.920 ;
  LAYER metal3 ;
  RECT 2938.580 1710.800 2942.120 1711.920 ;
  LAYER metal2 ;
  RECT 2938.580 1710.800 2942.120 1711.920 ;
  LAYER metal1 ;
  RECT 2938.580 1710.800 2942.120 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2929.900 1710.800 2933.440 1711.920 ;
  LAYER metal4 ;
  RECT 2929.900 1710.800 2933.440 1711.920 ;
  LAYER metal3 ;
  RECT 2929.900 1710.800 2933.440 1711.920 ;
  LAYER metal2 ;
  RECT 2929.900 1710.800 2933.440 1711.920 ;
  LAYER metal1 ;
  RECT 2929.900 1710.800 2933.440 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2921.220 1710.800 2924.760 1711.920 ;
  LAYER metal4 ;
  RECT 2921.220 1710.800 2924.760 1711.920 ;
  LAYER metal3 ;
  RECT 2921.220 1710.800 2924.760 1711.920 ;
  LAYER metal2 ;
  RECT 2921.220 1710.800 2924.760 1711.920 ;
  LAYER metal1 ;
  RECT 2921.220 1710.800 2924.760 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2877.820 1710.800 2881.360 1711.920 ;
  LAYER metal4 ;
  RECT 2877.820 1710.800 2881.360 1711.920 ;
  LAYER metal3 ;
  RECT 2877.820 1710.800 2881.360 1711.920 ;
  LAYER metal2 ;
  RECT 2877.820 1710.800 2881.360 1711.920 ;
  LAYER metal1 ;
  RECT 2877.820 1710.800 2881.360 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2869.140 1710.800 2872.680 1711.920 ;
  LAYER metal4 ;
  RECT 2869.140 1710.800 2872.680 1711.920 ;
  LAYER metal3 ;
  RECT 2869.140 1710.800 2872.680 1711.920 ;
  LAYER metal2 ;
  RECT 2869.140 1710.800 2872.680 1711.920 ;
  LAYER metal1 ;
  RECT 2869.140 1710.800 2872.680 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2860.460 1710.800 2864.000 1711.920 ;
  LAYER metal4 ;
  RECT 2860.460 1710.800 2864.000 1711.920 ;
  LAYER metal3 ;
  RECT 2860.460 1710.800 2864.000 1711.920 ;
  LAYER metal2 ;
  RECT 2860.460 1710.800 2864.000 1711.920 ;
  LAYER metal1 ;
  RECT 2860.460 1710.800 2864.000 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2851.780 1710.800 2855.320 1711.920 ;
  LAYER metal4 ;
  RECT 2851.780 1710.800 2855.320 1711.920 ;
  LAYER metal3 ;
  RECT 2851.780 1710.800 2855.320 1711.920 ;
  LAYER metal2 ;
  RECT 2851.780 1710.800 2855.320 1711.920 ;
  LAYER metal1 ;
  RECT 2851.780 1710.800 2855.320 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2843.100 1710.800 2846.640 1711.920 ;
  LAYER metal4 ;
  RECT 2843.100 1710.800 2846.640 1711.920 ;
  LAYER metal3 ;
  RECT 2843.100 1710.800 2846.640 1711.920 ;
  LAYER metal2 ;
  RECT 2843.100 1710.800 2846.640 1711.920 ;
  LAYER metal1 ;
  RECT 2843.100 1710.800 2846.640 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2834.420 1710.800 2837.960 1711.920 ;
  LAYER metal4 ;
  RECT 2834.420 1710.800 2837.960 1711.920 ;
  LAYER metal3 ;
  RECT 2834.420 1710.800 2837.960 1711.920 ;
  LAYER metal2 ;
  RECT 2834.420 1710.800 2837.960 1711.920 ;
  LAYER metal1 ;
  RECT 2834.420 1710.800 2837.960 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2791.020 1710.800 2794.560 1711.920 ;
  LAYER metal4 ;
  RECT 2791.020 1710.800 2794.560 1711.920 ;
  LAYER metal3 ;
  RECT 2791.020 1710.800 2794.560 1711.920 ;
  LAYER metal2 ;
  RECT 2791.020 1710.800 2794.560 1711.920 ;
  LAYER metal1 ;
  RECT 2791.020 1710.800 2794.560 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2782.340 1710.800 2785.880 1711.920 ;
  LAYER metal4 ;
  RECT 2782.340 1710.800 2785.880 1711.920 ;
  LAYER metal3 ;
  RECT 2782.340 1710.800 2785.880 1711.920 ;
  LAYER metal2 ;
  RECT 2782.340 1710.800 2785.880 1711.920 ;
  LAYER metal1 ;
  RECT 2782.340 1710.800 2785.880 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2769.320 1710.800 2772.860 1711.920 ;
  LAYER metal4 ;
  RECT 2769.320 1710.800 2772.860 1711.920 ;
  LAYER metal3 ;
  RECT 2769.320 1710.800 2772.860 1711.920 ;
  LAYER metal2 ;
  RECT 2769.320 1710.800 2772.860 1711.920 ;
  LAYER metal1 ;
  RECT 2769.320 1710.800 2772.860 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2755.680 1710.800 2759.220 1711.920 ;
  LAYER metal4 ;
  RECT 2755.680 1710.800 2759.220 1711.920 ;
  LAYER metal3 ;
  RECT 2755.680 1710.800 2759.220 1711.920 ;
  LAYER metal2 ;
  RECT 2755.680 1710.800 2759.220 1711.920 ;
  LAYER metal1 ;
  RECT 2755.680 1710.800 2759.220 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2742.040 1710.800 2745.580 1711.920 ;
  LAYER metal4 ;
  RECT 2742.040 1710.800 2745.580 1711.920 ;
  LAYER metal3 ;
  RECT 2742.040 1710.800 2745.580 1711.920 ;
  LAYER metal2 ;
  RECT 2742.040 1710.800 2745.580 1711.920 ;
  LAYER metal1 ;
  RECT 2742.040 1710.800 2745.580 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2727.780 1710.800 2731.320 1711.920 ;
  LAYER metal4 ;
  RECT 2727.780 1710.800 2731.320 1711.920 ;
  LAYER metal3 ;
  RECT 2727.780 1710.800 2731.320 1711.920 ;
  LAYER metal2 ;
  RECT 2727.780 1710.800 2731.320 1711.920 ;
  LAYER metal1 ;
  RECT 2727.780 1710.800 2731.320 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2684.380 1710.800 2687.920 1711.920 ;
  LAYER metal4 ;
  RECT 2684.380 1710.800 2687.920 1711.920 ;
  LAYER metal3 ;
  RECT 2684.380 1710.800 2687.920 1711.920 ;
  LAYER metal2 ;
  RECT 2684.380 1710.800 2687.920 1711.920 ;
  LAYER metal1 ;
  RECT 2684.380 1710.800 2687.920 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2675.700 1710.800 2679.240 1711.920 ;
  LAYER metal4 ;
  RECT 2675.700 1710.800 2679.240 1711.920 ;
  LAYER metal3 ;
  RECT 2675.700 1710.800 2679.240 1711.920 ;
  LAYER metal2 ;
  RECT 2675.700 1710.800 2679.240 1711.920 ;
  LAYER metal1 ;
  RECT 2675.700 1710.800 2679.240 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2667.020 1710.800 2670.560 1711.920 ;
  LAYER metal4 ;
  RECT 2667.020 1710.800 2670.560 1711.920 ;
  LAYER metal3 ;
  RECT 2667.020 1710.800 2670.560 1711.920 ;
  LAYER metal2 ;
  RECT 2667.020 1710.800 2670.560 1711.920 ;
  LAYER metal1 ;
  RECT 2667.020 1710.800 2670.560 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2658.340 1710.800 2661.880 1711.920 ;
  LAYER metal4 ;
  RECT 2658.340 1710.800 2661.880 1711.920 ;
  LAYER metal3 ;
  RECT 2658.340 1710.800 2661.880 1711.920 ;
  LAYER metal2 ;
  RECT 2658.340 1710.800 2661.880 1711.920 ;
  LAYER metal1 ;
  RECT 2658.340 1710.800 2661.880 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2649.660 1710.800 2653.200 1711.920 ;
  LAYER metal4 ;
  RECT 2649.660 1710.800 2653.200 1711.920 ;
  LAYER metal3 ;
  RECT 2649.660 1710.800 2653.200 1711.920 ;
  LAYER metal2 ;
  RECT 2649.660 1710.800 2653.200 1711.920 ;
  LAYER metal1 ;
  RECT 2649.660 1710.800 2653.200 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2640.980 1710.800 2644.520 1711.920 ;
  LAYER metal4 ;
  RECT 2640.980 1710.800 2644.520 1711.920 ;
  LAYER metal3 ;
  RECT 2640.980 1710.800 2644.520 1711.920 ;
  LAYER metal2 ;
  RECT 2640.980 1710.800 2644.520 1711.920 ;
  LAYER metal1 ;
  RECT 2640.980 1710.800 2644.520 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2597.580 1710.800 2601.120 1711.920 ;
  LAYER metal4 ;
  RECT 2597.580 1710.800 2601.120 1711.920 ;
  LAYER metal3 ;
  RECT 2597.580 1710.800 2601.120 1711.920 ;
  LAYER metal2 ;
  RECT 2597.580 1710.800 2601.120 1711.920 ;
  LAYER metal1 ;
  RECT 2597.580 1710.800 2601.120 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2588.900 1710.800 2592.440 1711.920 ;
  LAYER metal4 ;
  RECT 2588.900 1710.800 2592.440 1711.920 ;
  LAYER metal3 ;
  RECT 2588.900 1710.800 2592.440 1711.920 ;
  LAYER metal2 ;
  RECT 2588.900 1710.800 2592.440 1711.920 ;
  LAYER metal1 ;
  RECT 2588.900 1710.800 2592.440 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2580.220 1710.800 2583.760 1711.920 ;
  LAYER metal4 ;
  RECT 2580.220 1710.800 2583.760 1711.920 ;
  LAYER metal3 ;
  RECT 2580.220 1710.800 2583.760 1711.920 ;
  LAYER metal2 ;
  RECT 2580.220 1710.800 2583.760 1711.920 ;
  LAYER metal1 ;
  RECT 2580.220 1710.800 2583.760 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2571.540 1710.800 2575.080 1711.920 ;
  LAYER metal4 ;
  RECT 2571.540 1710.800 2575.080 1711.920 ;
  LAYER metal3 ;
  RECT 2571.540 1710.800 2575.080 1711.920 ;
  LAYER metal2 ;
  RECT 2571.540 1710.800 2575.080 1711.920 ;
  LAYER metal1 ;
  RECT 2571.540 1710.800 2575.080 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2562.860 1710.800 2566.400 1711.920 ;
  LAYER metal4 ;
  RECT 2562.860 1710.800 2566.400 1711.920 ;
  LAYER metal3 ;
  RECT 2562.860 1710.800 2566.400 1711.920 ;
  LAYER metal2 ;
  RECT 2562.860 1710.800 2566.400 1711.920 ;
  LAYER metal1 ;
  RECT 2562.860 1710.800 2566.400 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2554.180 1710.800 2557.720 1711.920 ;
  LAYER metal4 ;
  RECT 2554.180 1710.800 2557.720 1711.920 ;
  LAYER metal3 ;
  RECT 2554.180 1710.800 2557.720 1711.920 ;
  LAYER metal2 ;
  RECT 2554.180 1710.800 2557.720 1711.920 ;
  LAYER metal1 ;
  RECT 2554.180 1710.800 2557.720 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2510.780 1710.800 2514.320 1711.920 ;
  LAYER metal4 ;
  RECT 2510.780 1710.800 2514.320 1711.920 ;
  LAYER metal3 ;
  RECT 2510.780 1710.800 2514.320 1711.920 ;
  LAYER metal2 ;
  RECT 2510.780 1710.800 2514.320 1711.920 ;
  LAYER metal1 ;
  RECT 2510.780 1710.800 2514.320 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2502.100 1710.800 2505.640 1711.920 ;
  LAYER metal4 ;
  RECT 2502.100 1710.800 2505.640 1711.920 ;
  LAYER metal3 ;
  RECT 2502.100 1710.800 2505.640 1711.920 ;
  LAYER metal2 ;
  RECT 2502.100 1710.800 2505.640 1711.920 ;
  LAYER metal1 ;
  RECT 2502.100 1710.800 2505.640 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2493.420 1710.800 2496.960 1711.920 ;
  LAYER metal4 ;
  RECT 2493.420 1710.800 2496.960 1711.920 ;
  LAYER metal3 ;
  RECT 2493.420 1710.800 2496.960 1711.920 ;
  LAYER metal2 ;
  RECT 2493.420 1710.800 2496.960 1711.920 ;
  LAYER metal1 ;
  RECT 2493.420 1710.800 2496.960 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2484.740 1710.800 2488.280 1711.920 ;
  LAYER metal4 ;
  RECT 2484.740 1710.800 2488.280 1711.920 ;
  LAYER metal3 ;
  RECT 2484.740 1710.800 2488.280 1711.920 ;
  LAYER metal2 ;
  RECT 2484.740 1710.800 2488.280 1711.920 ;
  LAYER metal1 ;
  RECT 2484.740 1710.800 2488.280 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2476.060 1710.800 2479.600 1711.920 ;
  LAYER metal4 ;
  RECT 2476.060 1710.800 2479.600 1711.920 ;
  LAYER metal3 ;
  RECT 2476.060 1710.800 2479.600 1711.920 ;
  LAYER metal2 ;
  RECT 2476.060 1710.800 2479.600 1711.920 ;
  LAYER metal1 ;
  RECT 2476.060 1710.800 2479.600 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2467.380 1710.800 2470.920 1711.920 ;
  LAYER metal4 ;
  RECT 2467.380 1710.800 2470.920 1711.920 ;
  LAYER metal3 ;
  RECT 2467.380 1710.800 2470.920 1711.920 ;
  LAYER metal2 ;
  RECT 2467.380 1710.800 2470.920 1711.920 ;
  LAYER metal1 ;
  RECT 2467.380 1710.800 2470.920 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2423.980 1710.800 2427.520 1711.920 ;
  LAYER metal4 ;
  RECT 2423.980 1710.800 2427.520 1711.920 ;
  LAYER metal3 ;
  RECT 2423.980 1710.800 2427.520 1711.920 ;
  LAYER metal2 ;
  RECT 2423.980 1710.800 2427.520 1711.920 ;
  LAYER metal1 ;
  RECT 2423.980 1710.800 2427.520 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2415.300 1710.800 2418.840 1711.920 ;
  LAYER metal4 ;
  RECT 2415.300 1710.800 2418.840 1711.920 ;
  LAYER metal3 ;
  RECT 2415.300 1710.800 2418.840 1711.920 ;
  LAYER metal2 ;
  RECT 2415.300 1710.800 2418.840 1711.920 ;
  LAYER metal1 ;
  RECT 2415.300 1710.800 2418.840 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2406.620 1710.800 2410.160 1711.920 ;
  LAYER metal4 ;
  RECT 2406.620 1710.800 2410.160 1711.920 ;
  LAYER metal3 ;
  RECT 2406.620 1710.800 2410.160 1711.920 ;
  LAYER metal2 ;
  RECT 2406.620 1710.800 2410.160 1711.920 ;
  LAYER metal1 ;
  RECT 2406.620 1710.800 2410.160 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2397.940 1710.800 2401.480 1711.920 ;
  LAYER metal4 ;
  RECT 2397.940 1710.800 2401.480 1711.920 ;
  LAYER metal3 ;
  RECT 2397.940 1710.800 2401.480 1711.920 ;
  LAYER metal2 ;
  RECT 2397.940 1710.800 2401.480 1711.920 ;
  LAYER metal1 ;
  RECT 2397.940 1710.800 2401.480 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2389.260 1710.800 2392.800 1711.920 ;
  LAYER metal4 ;
  RECT 2389.260 1710.800 2392.800 1711.920 ;
  LAYER metal3 ;
  RECT 2389.260 1710.800 2392.800 1711.920 ;
  LAYER metal2 ;
  RECT 2389.260 1710.800 2392.800 1711.920 ;
  LAYER metal1 ;
  RECT 2389.260 1710.800 2392.800 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2380.580 1710.800 2384.120 1711.920 ;
  LAYER metal4 ;
  RECT 2380.580 1710.800 2384.120 1711.920 ;
  LAYER metal3 ;
  RECT 2380.580 1710.800 2384.120 1711.920 ;
  LAYER metal2 ;
  RECT 2380.580 1710.800 2384.120 1711.920 ;
  LAYER metal1 ;
  RECT 2380.580 1710.800 2384.120 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2327.880 1710.800 2331.420 1711.920 ;
  LAYER metal4 ;
  RECT 2327.880 1710.800 2331.420 1711.920 ;
  LAYER metal3 ;
  RECT 2327.880 1710.800 2331.420 1711.920 ;
  LAYER metal2 ;
  RECT 2327.880 1710.800 2331.420 1711.920 ;
  LAYER metal1 ;
  RECT 2327.880 1710.800 2331.420 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2314.240 1710.800 2317.780 1711.920 ;
  LAYER metal4 ;
  RECT 2314.240 1710.800 2317.780 1711.920 ;
  LAYER metal3 ;
  RECT 2314.240 1710.800 2317.780 1711.920 ;
  LAYER metal2 ;
  RECT 2314.240 1710.800 2317.780 1711.920 ;
  LAYER metal1 ;
  RECT 2314.240 1710.800 2317.780 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2299.980 1710.800 2303.520 1711.920 ;
  LAYER metal4 ;
  RECT 2299.980 1710.800 2303.520 1711.920 ;
  LAYER metal3 ;
  RECT 2299.980 1710.800 2303.520 1711.920 ;
  LAYER metal2 ;
  RECT 2299.980 1710.800 2303.520 1711.920 ;
  LAYER metal1 ;
  RECT 2299.980 1710.800 2303.520 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2291.300 1710.800 2294.840 1711.920 ;
  LAYER metal4 ;
  RECT 2291.300 1710.800 2294.840 1711.920 ;
  LAYER metal3 ;
  RECT 2291.300 1710.800 2294.840 1711.920 ;
  LAYER metal2 ;
  RECT 2291.300 1710.800 2294.840 1711.920 ;
  LAYER metal1 ;
  RECT 2291.300 1710.800 2294.840 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2282.620 1710.800 2286.160 1711.920 ;
  LAYER metal4 ;
  RECT 2282.620 1710.800 2286.160 1711.920 ;
  LAYER metal3 ;
  RECT 2282.620 1710.800 2286.160 1711.920 ;
  LAYER metal2 ;
  RECT 2282.620 1710.800 2286.160 1711.920 ;
  LAYER metal1 ;
  RECT 2282.620 1710.800 2286.160 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2273.940 1710.800 2277.480 1711.920 ;
  LAYER metal4 ;
  RECT 2273.940 1710.800 2277.480 1711.920 ;
  LAYER metal3 ;
  RECT 2273.940 1710.800 2277.480 1711.920 ;
  LAYER metal2 ;
  RECT 2273.940 1710.800 2277.480 1711.920 ;
  LAYER metal1 ;
  RECT 2273.940 1710.800 2277.480 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2230.540 1710.800 2234.080 1711.920 ;
  LAYER metal4 ;
  RECT 2230.540 1710.800 2234.080 1711.920 ;
  LAYER metal3 ;
  RECT 2230.540 1710.800 2234.080 1711.920 ;
  LAYER metal2 ;
  RECT 2230.540 1710.800 2234.080 1711.920 ;
  LAYER metal1 ;
  RECT 2230.540 1710.800 2234.080 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2221.860 1710.800 2225.400 1711.920 ;
  LAYER metal4 ;
  RECT 2221.860 1710.800 2225.400 1711.920 ;
  LAYER metal3 ;
  RECT 2221.860 1710.800 2225.400 1711.920 ;
  LAYER metal2 ;
  RECT 2221.860 1710.800 2225.400 1711.920 ;
  LAYER metal1 ;
  RECT 2221.860 1710.800 2225.400 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2213.180 1710.800 2216.720 1711.920 ;
  LAYER metal4 ;
  RECT 2213.180 1710.800 2216.720 1711.920 ;
  LAYER metal3 ;
  RECT 2213.180 1710.800 2216.720 1711.920 ;
  LAYER metal2 ;
  RECT 2213.180 1710.800 2216.720 1711.920 ;
  LAYER metal1 ;
  RECT 2213.180 1710.800 2216.720 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2204.500 1710.800 2208.040 1711.920 ;
  LAYER metal4 ;
  RECT 2204.500 1710.800 2208.040 1711.920 ;
  LAYER metal3 ;
  RECT 2204.500 1710.800 2208.040 1711.920 ;
  LAYER metal2 ;
  RECT 2204.500 1710.800 2208.040 1711.920 ;
  LAYER metal1 ;
  RECT 2204.500 1710.800 2208.040 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2195.820 1710.800 2199.360 1711.920 ;
  LAYER metal4 ;
  RECT 2195.820 1710.800 2199.360 1711.920 ;
  LAYER metal3 ;
  RECT 2195.820 1710.800 2199.360 1711.920 ;
  LAYER metal2 ;
  RECT 2195.820 1710.800 2199.360 1711.920 ;
  LAYER metal1 ;
  RECT 2195.820 1710.800 2199.360 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2187.140 1710.800 2190.680 1711.920 ;
  LAYER metal4 ;
  RECT 2187.140 1710.800 2190.680 1711.920 ;
  LAYER metal3 ;
  RECT 2187.140 1710.800 2190.680 1711.920 ;
  LAYER metal2 ;
  RECT 2187.140 1710.800 2190.680 1711.920 ;
  LAYER metal1 ;
  RECT 2187.140 1710.800 2190.680 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2143.740 1710.800 2147.280 1711.920 ;
  LAYER metal4 ;
  RECT 2143.740 1710.800 2147.280 1711.920 ;
  LAYER metal3 ;
  RECT 2143.740 1710.800 2147.280 1711.920 ;
  LAYER metal2 ;
  RECT 2143.740 1710.800 2147.280 1711.920 ;
  LAYER metal1 ;
  RECT 2143.740 1710.800 2147.280 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2135.060 1710.800 2138.600 1711.920 ;
  LAYER metal4 ;
  RECT 2135.060 1710.800 2138.600 1711.920 ;
  LAYER metal3 ;
  RECT 2135.060 1710.800 2138.600 1711.920 ;
  LAYER metal2 ;
  RECT 2135.060 1710.800 2138.600 1711.920 ;
  LAYER metal1 ;
  RECT 2135.060 1710.800 2138.600 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2126.380 1710.800 2129.920 1711.920 ;
  LAYER metal4 ;
  RECT 2126.380 1710.800 2129.920 1711.920 ;
  LAYER metal3 ;
  RECT 2126.380 1710.800 2129.920 1711.920 ;
  LAYER metal2 ;
  RECT 2126.380 1710.800 2129.920 1711.920 ;
  LAYER metal1 ;
  RECT 2126.380 1710.800 2129.920 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2117.700 1710.800 2121.240 1711.920 ;
  LAYER metal4 ;
  RECT 2117.700 1710.800 2121.240 1711.920 ;
  LAYER metal3 ;
  RECT 2117.700 1710.800 2121.240 1711.920 ;
  LAYER metal2 ;
  RECT 2117.700 1710.800 2121.240 1711.920 ;
  LAYER metal1 ;
  RECT 2117.700 1710.800 2121.240 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2109.020 1710.800 2112.560 1711.920 ;
  LAYER metal4 ;
  RECT 2109.020 1710.800 2112.560 1711.920 ;
  LAYER metal3 ;
  RECT 2109.020 1710.800 2112.560 1711.920 ;
  LAYER metal2 ;
  RECT 2109.020 1710.800 2112.560 1711.920 ;
  LAYER metal1 ;
  RECT 2109.020 1710.800 2112.560 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2100.340 1710.800 2103.880 1711.920 ;
  LAYER metal4 ;
  RECT 2100.340 1710.800 2103.880 1711.920 ;
  LAYER metal3 ;
  RECT 2100.340 1710.800 2103.880 1711.920 ;
  LAYER metal2 ;
  RECT 2100.340 1710.800 2103.880 1711.920 ;
  LAYER metal1 ;
  RECT 2100.340 1710.800 2103.880 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2056.940 1710.800 2060.480 1711.920 ;
  LAYER metal4 ;
  RECT 2056.940 1710.800 2060.480 1711.920 ;
  LAYER metal3 ;
  RECT 2056.940 1710.800 2060.480 1711.920 ;
  LAYER metal2 ;
  RECT 2056.940 1710.800 2060.480 1711.920 ;
  LAYER metal1 ;
  RECT 2056.940 1710.800 2060.480 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2048.260 1710.800 2051.800 1711.920 ;
  LAYER metal4 ;
  RECT 2048.260 1710.800 2051.800 1711.920 ;
  LAYER metal3 ;
  RECT 2048.260 1710.800 2051.800 1711.920 ;
  LAYER metal2 ;
  RECT 2048.260 1710.800 2051.800 1711.920 ;
  LAYER metal1 ;
  RECT 2048.260 1710.800 2051.800 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2039.580 1710.800 2043.120 1711.920 ;
  LAYER metal4 ;
  RECT 2039.580 1710.800 2043.120 1711.920 ;
  LAYER metal3 ;
  RECT 2039.580 1710.800 2043.120 1711.920 ;
  LAYER metal2 ;
  RECT 2039.580 1710.800 2043.120 1711.920 ;
  LAYER metal1 ;
  RECT 2039.580 1710.800 2043.120 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2030.900 1710.800 2034.440 1711.920 ;
  LAYER metal4 ;
  RECT 2030.900 1710.800 2034.440 1711.920 ;
  LAYER metal3 ;
  RECT 2030.900 1710.800 2034.440 1711.920 ;
  LAYER metal2 ;
  RECT 2030.900 1710.800 2034.440 1711.920 ;
  LAYER metal1 ;
  RECT 2030.900 1710.800 2034.440 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2022.220 1710.800 2025.760 1711.920 ;
  LAYER metal4 ;
  RECT 2022.220 1710.800 2025.760 1711.920 ;
  LAYER metal3 ;
  RECT 2022.220 1710.800 2025.760 1711.920 ;
  LAYER metal2 ;
  RECT 2022.220 1710.800 2025.760 1711.920 ;
  LAYER metal1 ;
  RECT 2022.220 1710.800 2025.760 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2013.540 1710.800 2017.080 1711.920 ;
  LAYER metal4 ;
  RECT 2013.540 1710.800 2017.080 1711.920 ;
  LAYER metal3 ;
  RECT 2013.540 1710.800 2017.080 1711.920 ;
  LAYER metal2 ;
  RECT 2013.540 1710.800 2017.080 1711.920 ;
  LAYER metal1 ;
  RECT 2013.540 1710.800 2017.080 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1970.140 1710.800 1973.680 1711.920 ;
  LAYER metal4 ;
  RECT 1970.140 1710.800 1973.680 1711.920 ;
  LAYER metal3 ;
  RECT 1970.140 1710.800 1973.680 1711.920 ;
  LAYER metal2 ;
  RECT 1970.140 1710.800 1973.680 1711.920 ;
  LAYER metal1 ;
  RECT 1970.140 1710.800 1973.680 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1961.460 1710.800 1965.000 1711.920 ;
  LAYER metal4 ;
  RECT 1961.460 1710.800 1965.000 1711.920 ;
  LAYER metal3 ;
  RECT 1961.460 1710.800 1965.000 1711.920 ;
  LAYER metal2 ;
  RECT 1961.460 1710.800 1965.000 1711.920 ;
  LAYER metal1 ;
  RECT 1961.460 1710.800 1965.000 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1952.780 1710.800 1956.320 1711.920 ;
  LAYER metal4 ;
  RECT 1952.780 1710.800 1956.320 1711.920 ;
  LAYER metal3 ;
  RECT 1952.780 1710.800 1956.320 1711.920 ;
  LAYER metal2 ;
  RECT 1952.780 1710.800 1956.320 1711.920 ;
  LAYER metal1 ;
  RECT 1952.780 1710.800 1956.320 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1944.100 1710.800 1947.640 1711.920 ;
  LAYER metal4 ;
  RECT 1944.100 1710.800 1947.640 1711.920 ;
  LAYER metal3 ;
  RECT 1944.100 1710.800 1947.640 1711.920 ;
  LAYER metal2 ;
  RECT 1944.100 1710.800 1947.640 1711.920 ;
  LAYER metal1 ;
  RECT 1944.100 1710.800 1947.640 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1935.420 1710.800 1938.960 1711.920 ;
  LAYER metal4 ;
  RECT 1935.420 1710.800 1938.960 1711.920 ;
  LAYER metal3 ;
  RECT 1935.420 1710.800 1938.960 1711.920 ;
  LAYER metal2 ;
  RECT 1935.420 1710.800 1938.960 1711.920 ;
  LAYER metal1 ;
  RECT 1935.420 1710.800 1938.960 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1926.740 1710.800 1930.280 1711.920 ;
  LAYER metal4 ;
  RECT 1926.740 1710.800 1930.280 1711.920 ;
  LAYER metal3 ;
  RECT 1926.740 1710.800 1930.280 1711.920 ;
  LAYER metal2 ;
  RECT 1926.740 1710.800 1930.280 1711.920 ;
  LAYER metal1 ;
  RECT 1926.740 1710.800 1930.280 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1863.500 1710.800 1867.040 1711.920 ;
  LAYER metal4 ;
  RECT 1863.500 1710.800 1867.040 1711.920 ;
  LAYER metal3 ;
  RECT 1863.500 1710.800 1867.040 1711.920 ;
  LAYER metal2 ;
  RECT 1863.500 1710.800 1867.040 1711.920 ;
  LAYER metal1 ;
  RECT 1863.500 1710.800 1867.040 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1854.820 1710.800 1858.360 1711.920 ;
  LAYER metal4 ;
  RECT 1854.820 1710.800 1858.360 1711.920 ;
  LAYER metal3 ;
  RECT 1854.820 1710.800 1858.360 1711.920 ;
  LAYER metal2 ;
  RECT 1854.820 1710.800 1858.360 1711.920 ;
  LAYER metal1 ;
  RECT 1854.820 1710.800 1858.360 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1813.280 1710.800 1816.820 1711.920 ;
  LAYER metal4 ;
  RECT 1813.280 1710.800 1816.820 1711.920 ;
  LAYER metal3 ;
  RECT 1813.280 1710.800 1816.820 1711.920 ;
  LAYER metal2 ;
  RECT 1813.280 1710.800 1816.820 1711.920 ;
  LAYER metal1 ;
  RECT 1813.280 1710.800 1816.820 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1789.100 1710.800 1792.640 1711.920 ;
  LAYER metal4 ;
  RECT 1789.100 1710.800 1792.640 1711.920 ;
  LAYER metal3 ;
  RECT 1789.100 1710.800 1792.640 1711.920 ;
  LAYER metal2 ;
  RECT 1789.100 1710.800 1792.640 1711.920 ;
  LAYER metal1 ;
  RECT 1789.100 1710.800 1792.640 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1764.300 1710.800 1767.840 1711.920 ;
  LAYER metal4 ;
  RECT 1764.300 1710.800 1767.840 1711.920 ;
  LAYER metal3 ;
  RECT 1764.300 1710.800 1767.840 1711.920 ;
  LAYER metal2 ;
  RECT 1764.300 1710.800 1767.840 1711.920 ;
  LAYER metal1 ;
  RECT 1764.300 1710.800 1767.840 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1738.260 1710.800 1741.800 1711.920 ;
  LAYER metal4 ;
  RECT 1738.260 1710.800 1741.800 1711.920 ;
  LAYER metal3 ;
  RECT 1738.260 1710.800 1741.800 1711.920 ;
  LAYER metal2 ;
  RECT 1738.260 1710.800 1741.800 1711.920 ;
  LAYER metal1 ;
  RECT 1738.260 1710.800 1741.800 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1694.860 1710.800 1698.400 1711.920 ;
  LAYER metal4 ;
  RECT 1694.860 1710.800 1698.400 1711.920 ;
  LAYER metal3 ;
  RECT 1694.860 1710.800 1698.400 1711.920 ;
  LAYER metal2 ;
  RECT 1694.860 1710.800 1698.400 1711.920 ;
  LAYER metal1 ;
  RECT 1694.860 1710.800 1698.400 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1686.180 1710.800 1689.720 1711.920 ;
  LAYER metal4 ;
  RECT 1686.180 1710.800 1689.720 1711.920 ;
  LAYER metal3 ;
  RECT 1686.180 1710.800 1689.720 1711.920 ;
  LAYER metal2 ;
  RECT 1686.180 1710.800 1689.720 1711.920 ;
  LAYER metal1 ;
  RECT 1686.180 1710.800 1689.720 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1677.500 1710.800 1681.040 1711.920 ;
  LAYER metal4 ;
  RECT 1677.500 1710.800 1681.040 1711.920 ;
  LAYER metal3 ;
  RECT 1677.500 1710.800 1681.040 1711.920 ;
  LAYER metal2 ;
  RECT 1677.500 1710.800 1681.040 1711.920 ;
  LAYER metal1 ;
  RECT 1677.500 1710.800 1681.040 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1668.820 1710.800 1672.360 1711.920 ;
  LAYER metal4 ;
  RECT 1668.820 1710.800 1672.360 1711.920 ;
  LAYER metal3 ;
  RECT 1668.820 1710.800 1672.360 1711.920 ;
  LAYER metal2 ;
  RECT 1668.820 1710.800 1672.360 1711.920 ;
  LAYER metal1 ;
  RECT 1668.820 1710.800 1672.360 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1660.140 1710.800 1663.680 1711.920 ;
  LAYER metal4 ;
  RECT 1660.140 1710.800 1663.680 1711.920 ;
  LAYER metal3 ;
  RECT 1660.140 1710.800 1663.680 1711.920 ;
  LAYER metal2 ;
  RECT 1660.140 1710.800 1663.680 1711.920 ;
  LAYER metal1 ;
  RECT 1660.140 1710.800 1663.680 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1651.460 1710.800 1655.000 1711.920 ;
  LAYER metal4 ;
  RECT 1651.460 1710.800 1655.000 1711.920 ;
  LAYER metal3 ;
  RECT 1651.460 1710.800 1655.000 1711.920 ;
  LAYER metal2 ;
  RECT 1651.460 1710.800 1655.000 1711.920 ;
  LAYER metal1 ;
  RECT 1651.460 1710.800 1655.000 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1608.060 1710.800 1611.600 1711.920 ;
  LAYER metal4 ;
  RECT 1608.060 1710.800 1611.600 1711.920 ;
  LAYER metal3 ;
  RECT 1608.060 1710.800 1611.600 1711.920 ;
  LAYER metal2 ;
  RECT 1608.060 1710.800 1611.600 1711.920 ;
  LAYER metal1 ;
  RECT 1608.060 1710.800 1611.600 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1599.380 1710.800 1602.920 1711.920 ;
  LAYER metal4 ;
  RECT 1599.380 1710.800 1602.920 1711.920 ;
  LAYER metal3 ;
  RECT 1599.380 1710.800 1602.920 1711.920 ;
  LAYER metal2 ;
  RECT 1599.380 1710.800 1602.920 1711.920 ;
  LAYER metal1 ;
  RECT 1599.380 1710.800 1602.920 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1590.700 1710.800 1594.240 1711.920 ;
  LAYER metal4 ;
  RECT 1590.700 1710.800 1594.240 1711.920 ;
  LAYER metal3 ;
  RECT 1590.700 1710.800 1594.240 1711.920 ;
  LAYER metal2 ;
  RECT 1590.700 1710.800 1594.240 1711.920 ;
  LAYER metal1 ;
  RECT 1590.700 1710.800 1594.240 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1582.020 1710.800 1585.560 1711.920 ;
  LAYER metal4 ;
  RECT 1582.020 1710.800 1585.560 1711.920 ;
  LAYER metal3 ;
  RECT 1582.020 1710.800 1585.560 1711.920 ;
  LAYER metal2 ;
  RECT 1582.020 1710.800 1585.560 1711.920 ;
  LAYER metal1 ;
  RECT 1582.020 1710.800 1585.560 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1573.340 1710.800 1576.880 1711.920 ;
  LAYER metal4 ;
  RECT 1573.340 1710.800 1576.880 1711.920 ;
  LAYER metal3 ;
  RECT 1573.340 1710.800 1576.880 1711.920 ;
  LAYER metal2 ;
  RECT 1573.340 1710.800 1576.880 1711.920 ;
  LAYER metal1 ;
  RECT 1573.340 1710.800 1576.880 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1564.660 1710.800 1568.200 1711.920 ;
  LAYER metal4 ;
  RECT 1564.660 1710.800 1568.200 1711.920 ;
  LAYER metal3 ;
  RECT 1564.660 1710.800 1568.200 1711.920 ;
  LAYER metal2 ;
  RECT 1564.660 1710.800 1568.200 1711.920 ;
  LAYER metal1 ;
  RECT 1564.660 1710.800 1568.200 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1521.260 1710.800 1524.800 1711.920 ;
  LAYER metal4 ;
  RECT 1521.260 1710.800 1524.800 1711.920 ;
  LAYER metal3 ;
  RECT 1521.260 1710.800 1524.800 1711.920 ;
  LAYER metal2 ;
  RECT 1521.260 1710.800 1524.800 1711.920 ;
  LAYER metal1 ;
  RECT 1521.260 1710.800 1524.800 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1512.580 1710.800 1516.120 1711.920 ;
  LAYER metal4 ;
  RECT 1512.580 1710.800 1516.120 1711.920 ;
  LAYER metal3 ;
  RECT 1512.580 1710.800 1516.120 1711.920 ;
  LAYER metal2 ;
  RECT 1512.580 1710.800 1516.120 1711.920 ;
  LAYER metal1 ;
  RECT 1512.580 1710.800 1516.120 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1503.900 1710.800 1507.440 1711.920 ;
  LAYER metal4 ;
  RECT 1503.900 1710.800 1507.440 1711.920 ;
  LAYER metal3 ;
  RECT 1503.900 1710.800 1507.440 1711.920 ;
  LAYER metal2 ;
  RECT 1503.900 1710.800 1507.440 1711.920 ;
  LAYER metal1 ;
  RECT 1503.900 1710.800 1507.440 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1495.220 1710.800 1498.760 1711.920 ;
  LAYER metal4 ;
  RECT 1495.220 1710.800 1498.760 1711.920 ;
  LAYER metal3 ;
  RECT 1495.220 1710.800 1498.760 1711.920 ;
  LAYER metal2 ;
  RECT 1495.220 1710.800 1498.760 1711.920 ;
  LAYER metal1 ;
  RECT 1495.220 1710.800 1498.760 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1486.540 1710.800 1490.080 1711.920 ;
  LAYER metal4 ;
  RECT 1486.540 1710.800 1490.080 1711.920 ;
  LAYER metal3 ;
  RECT 1486.540 1710.800 1490.080 1711.920 ;
  LAYER metal2 ;
  RECT 1486.540 1710.800 1490.080 1711.920 ;
  LAYER metal1 ;
  RECT 1486.540 1710.800 1490.080 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1477.860 1710.800 1481.400 1711.920 ;
  LAYER metal4 ;
  RECT 1477.860 1710.800 1481.400 1711.920 ;
  LAYER metal3 ;
  RECT 1477.860 1710.800 1481.400 1711.920 ;
  LAYER metal2 ;
  RECT 1477.860 1710.800 1481.400 1711.920 ;
  LAYER metal1 ;
  RECT 1477.860 1710.800 1481.400 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1434.460 1710.800 1438.000 1711.920 ;
  LAYER metal4 ;
  RECT 1434.460 1710.800 1438.000 1711.920 ;
  LAYER metal3 ;
  RECT 1434.460 1710.800 1438.000 1711.920 ;
  LAYER metal2 ;
  RECT 1434.460 1710.800 1438.000 1711.920 ;
  LAYER metal1 ;
  RECT 1434.460 1710.800 1438.000 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1425.780 1710.800 1429.320 1711.920 ;
  LAYER metal4 ;
  RECT 1425.780 1710.800 1429.320 1711.920 ;
  LAYER metal3 ;
  RECT 1425.780 1710.800 1429.320 1711.920 ;
  LAYER metal2 ;
  RECT 1425.780 1710.800 1429.320 1711.920 ;
  LAYER metal1 ;
  RECT 1425.780 1710.800 1429.320 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1417.100 1710.800 1420.640 1711.920 ;
  LAYER metal4 ;
  RECT 1417.100 1710.800 1420.640 1711.920 ;
  LAYER metal3 ;
  RECT 1417.100 1710.800 1420.640 1711.920 ;
  LAYER metal2 ;
  RECT 1417.100 1710.800 1420.640 1711.920 ;
  LAYER metal1 ;
  RECT 1417.100 1710.800 1420.640 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1408.420 1710.800 1411.960 1711.920 ;
  LAYER metal4 ;
  RECT 1408.420 1710.800 1411.960 1711.920 ;
  LAYER metal3 ;
  RECT 1408.420 1710.800 1411.960 1711.920 ;
  LAYER metal2 ;
  RECT 1408.420 1710.800 1411.960 1711.920 ;
  LAYER metal1 ;
  RECT 1408.420 1710.800 1411.960 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1399.740 1710.800 1403.280 1711.920 ;
  LAYER metal4 ;
  RECT 1399.740 1710.800 1403.280 1711.920 ;
  LAYER metal3 ;
  RECT 1399.740 1710.800 1403.280 1711.920 ;
  LAYER metal2 ;
  RECT 1399.740 1710.800 1403.280 1711.920 ;
  LAYER metal1 ;
  RECT 1399.740 1710.800 1403.280 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1391.060 1710.800 1394.600 1711.920 ;
  LAYER metal4 ;
  RECT 1391.060 1710.800 1394.600 1711.920 ;
  LAYER metal3 ;
  RECT 1391.060 1710.800 1394.600 1711.920 ;
  LAYER metal2 ;
  RECT 1391.060 1710.800 1394.600 1711.920 ;
  LAYER metal1 ;
  RECT 1391.060 1710.800 1394.600 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1343.320 1710.800 1346.860 1711.920 ;
  LAYER metal4 ;
  RECT 1343.320 1710.800 1346.860 1711.920 ;
  LAYER metal3 ;
  RECT 1343.320 1710.800 1346.860 1711.920 ;
  LAYER metal2 ;
  RECT 1343.320 1710.800 1346.860 1711.920 ;
  LAYER metal1 ;
  RECT 1343.320 1710.800 1346.860 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1329.680 1710.800 1333.220 1711.920 ;
  LAYER metal4 ;
  RECT 1329.680 1710.800 1333.220 1711.920 ;
  LAYER metal3 ;
  RECT 1329.680 1710.800 1333.220 1711.920 ;
  LAYER metal2 ;
  RECT 1329.680 1710.800 1333.220 1711.920 ;
  LAYER metal1 ;
  RECT 1329.680 1710.800 1333.220 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1316.040 1710.800 1319.580 1711.920 ;
  LAYER metal4 ;
  RECT 1316.040 1710.800 1319.580 1711.920 ;
  LAYER metal3 ;
  RECT 1316.040 1710.800 1319.580 1711.920 ;
  LAYER metal2 ;
  RECT 1316.040 1710.800 1319.580 1711.920 ;
  LAYER metal1 ;
  RECT 1316.040 1710.800 1319.580 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1301.780 1710.800 1305.320 1711.920 ;
  LAYER metal4 ;
  RECT 1301.780 1710.800 1305.320 1711.920 ;
  LAYER metal3 ;
  RECT 1301.780 1710.800 1305.320 1711.920 ;
  LAYER metal2 ;
  RECT 1301.780 1710.800 1305.320 1711.920 ;
  LAYER metal1 ;
  RECT 1301.780 1710.800 1305.320 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1293.100 1710.800 1296.640 1711.920 ;
  LAYER metal4 ;
  RECT 1293.100 1710.800 1296.640 1711.920 ;
  LAYER metal3 ;
  RECT 1293.100 1710.800 1296.640 1711.920 ;
  LAYER metal2 ;
  RECT 1293.100 1710.800 1296.640 1711.920 ;
  LAYER metal1 ;
  RECT 1293.100 1710.800 1296.640 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1284.420 1710.800 1287.960 1711.920 ;
  LAYER metal4 ;
  RECT 1284.420 1710.800 1287.960 1711.920 ;
  LAYER metal3 ;
  RECT 1284.420 1710.800 1287.960 1711.920 ;
  LAYER metal2 ;
  RECT 1284.420 1710.800 1287.960 1711.920 ;
  LAYER metal1 ;
  RECT 1284.420 1710.800 1287.960 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1241.020 1710.800 1244.560 1711.920 ;
  LAYER metal4 ;
  RECT 1241.020 1710.800 1244.560 1711.920 ;
  LAYER metal3 ;
  RECT 1241.020 1710.800 1244.560 1711.920 ;
  LAYER metal2 ;
  RECT 1241.020 1710.800 1244.560 1711.920 ;
  LAYER metal1 ;
  RECT 1241.020 1710.800 1244.560 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1232.340 1710.800 1235.880 1711.920 ;
  LAYER metal4 ;
  RECT 1232.340 1710.800 1235.880 1711.920 ;
  LAYER metal3 ;
  RECT 1232.340 1710.800 1235.880 1711.920 ;
  LAYER metal2 ;
  RECT 1232.340 1710.800 1235.880 1711.920 ;
  LAYER metal1 ;
  RECT 1232.340 1710.800 1235.880 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1223.660 1710.800 1227.200 1711.920 ;
  LAYER metal4 ;
  RECT 1223.660 1710.800 1227.200 1711.920 ;
  LAYER metal3 ;
  RECT 1223.660 1710.800 1227.200 1711.920 ;
  LAYER metal2 ;
  RECT 1223.660 1710.800 1227.200 1711.920 ;
  LAYER metal1 ;
  RECT 1223.660 1710.800 1227.200 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1214.980 1710.800 1218.520 1711.920 ;
  LAYER metal4 ;
  RECT 1214.980 1710.800 1218.520 1711.920 ;
  LAYER metal3 ;
  RECT 1214.980 1710.800 1218.520 1711.920 ;
  LAYER metal2 ;
  RECT 1214.980 1710.800 1218.520 1711.920 ;
  LAYER metal1 ;
  RECT 1214.980 1710.800 1218.520 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1206.300 1710.800 1209.840 1711.920 ;
  LAYER metal4 ;
  RECT 1206.300 1710.800 1209.840 1711.920 ;
  LAYER metal3 ;
  RECT 1206.300 1710.800 1209.840 1711.920 ;
  LAYER metal2 ;
  RECT 1206.300 1710.800 1209.840 1711.920 ;
  LAYER metal1 ;
  RECT 1206.300 1710.800 1209.840 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1197.620 1710.800 1201.160 1711.920 ;
  LAYER metal4 ;
  RECT 1197.620 1710.800 1201.160 1711.920 ;
  LAYER metal3 ;
  RECT 1197.620 1710.800 1201.160 1711.920 ;
  LAYER metal2 ;
  RECT 1197.620 1710.800 1201.160 1711.920 ;
  LAYER metal1 ;
  RECT 1197.620 1710.800 1201.160 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1154.220 1710.800 1157.760 1711.920 ;
  LAYER metal4 ;
  RECT 1154.220 1710.800 1157.760 1711.920 ;
  LAYER metal3 ;
  RECT 1154.220 1710.800 1157.760 1711.920 ;
  LAYER metal2 ;
  RECT 1154.220 1710.800 1157.760 1711.920 ;
  LAYER metal1 ;
  RECT 1154.220 1710.800 1157.760 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1145.540 1710.800 1149.080 1711.920 ;
  LAYER metal4 ;
  RECT 1145.540 1710.800 1149.080 1711.920 ;
  LAYER metal3 ;
  RECT 1145.540 1710.800 1149.080 1711.920 ;
  LAYER metal2 ;
  RECT 1145.540 1710.800 1149.080 1711.920 ;
  LAYER metal1 ;
  RECT 1145.540 1710.800 1149.080 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1136.860 1710.800 1140.400 1711.920 ;
  LAYER metal4 ;
  RECT 1136.860 1710.800 1140.400 1711.920 ;
  LAYER metal3 ;
  RECT 1136.860 1710.800 1140.400 1711.920 ;
  LAYER metal2 ;
  RECT 1136.860 1710.800 1140.400 1711.920 ;
  LAYER metal1 ;
  RECT 1136.860 1710.800 1140.400 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1128.180 1710.800 1131.720 1711.920 ;
  LAYER metal4 ;
  RECT 1128.180 1710.800 1131.720 1711.920 ;
  LAYER metal3 ;
  RECT 1128.180 1710.800 1131.720 1711.920 ;
  LAYER metal2 ;
  RECT 1128.180 1710.800 1131.720 1711.920 ;
  LAYER metal1 ;
  RECT 1128.180 1710.800 1131.720 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1119.500 1710.800 1123.040 1711.920 ;
  LAYER metal4 ;
  RECT 1119.500 1710.800 1123.040 1711.920 ;
  LAYER metal3 ;
  RECT 1119.500 1710.800 1123.040 1711.920 ;
  LAYER metal2 ;
  RECT 1119.500 1710.800 1123.040 1711.920 ;
  LAYER metal1 ;
  RECT 1119.500 1710.800 1123.040 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1110.820 1710.800 1114.360 1711.920 ;
  LAYER metal4 ;
  RECT 1110.820 1710.800 1114.360 1711.920 ;
  LAYER metal3 ;
  RECT 1110.820 1710.800 1114.360 1711.920 ;
  LAYER metal2 ;
  RECT 1110.820 1710.800 1114.360 1711.920 ;
  LAYER metal1 ;
  RECT 1110.820 1710.800 1114.360 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1067.420 1710.800 1070.960 1711.920 ;
  LAYER metal4 ;
  RECT 1067.420 1710.800 1070.960 1711.920 ;
  LAYER metal3 ;
  RECT 1067.420 1710.800 1070.960 1711.920 ;
  LAYER metal2 ;
  RECT 1067.420 1710.800 1070.960 1711.920 ;
  LAYER metal1 ;
  RECT 1067.420 1710.800 1070.960 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1058.740 1710.800 1062.280 1711.920 ;
  LAYER metal4 ;
  RECT 1058.740 1710.800 1062.280 1711.920 ;
  LAYER metal3 ;
  RECT 1058.740 1710.800 1062.280 1711.920 ;
  LAYER metal2 ;
  RECT 1058.740 1710.800 1062.280 1711.920 ;
  LAYER metal1 ;
  RECT 1058.740 1710.800 1062.280 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1050.060 1710.800 1053.600 1711.920 ;
  LAYER metal4 ;
  RECT 1050.060 1710.800 1053.600 1711.920 ;
  LAYER metal3 ;
  RECT 1050.060 1710.800 1053.600 1711.920 ;
  LAYER metal2 ;
  RECT 1050.060 1710.800 1053.600 1711.920 ;
  LAYER metal1 ;
  RECT 1050.060 1710.800 1053.600 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1041.380 1710.800 1044.920 1711.920 ;
  LAYER metal4 ;
  RECT 1041.380 1710.800 1044.920 1711.920 ;
  LAYER metal3 ;
  RECT 1041.380 1710.800 1044.920 1711.920 ;
  LAYER metal2 ;
  RECT 1041.380 1710.800 1044.920 1711.920 ;
  LAYER metal1 ;
  RECT 1041.380 1710.800 1044.920 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1032.700 1710.800 1036.240 1711.920 ;
  LAYER metal4 ;
  RECT 1032.700 1710.800 1036.240 1711.920 ;
  LAYER metal3 ;
  RECT 1032.700 1710.800 1036.240 1711.920 ;
  LAYER metal2 ;
  RECT 1032.700 1710.800 1036.240 1711.920 ;
  LAYER metal1 ;
  RECT 1032.700 1710.800 1036.240 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1024.020 1710.800 1027.560 1711.920 ;
  LAYER metal4 ;
  RECT 1024.020 1710.800 1027.560 1711.920 ;
  LAYER metal3 ;
  RECT 1024.020 1710.800 1027.560 1711.920 ;
  LAYER metal2 ;
  RECT 1024.020 1710.800 1027.560 1711.920 ;
  LAYER metal1 ;
  RECT 1024.020 1710.800 1027.560 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 980.620 1710.800 984.160 1711.920 ;
  LAYER metal4 ;
  RECT 980.620 1710.800 984.160 1711.920 ;
  LAYER metal3 ;
  RECT 980.620 1710.800 984.160 1711.920 ;
  LAYER metal2 ;
  RECT 980.620 1710.800 984.160 1711.920 ;
  LAYER metal1 ;
  RECT 980.620 1710.800 984.160 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 971.940 1710.800 975.480 1711.920 ;
  LAYER metal4 ;
  RECT 971.940 1710.800 975.480 1711.920 ;
  LAYER metal3 ;
  RECT 971.940 1710.800 975.480 1711.920 ;
  LAYER metal2 ;
  RECT 971.940 1710.800 975.480 1711.920 ;
  LAYER metal1 ;
  RECT 971.940 1710.800 975.480 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 963.260 1710.800 966.800 1711.920 ;
  LAYER metal4 ;
  RECT 963.260 1710.800 966.800 1711.920 ;
  LAYER metal3 ;
  RECT 963.260 1710.800 966.800 1711.920 ;
  LAYER metal2 ;
  RECT 963.260 1710.800 966.800 1711.920 ;
  LAYER metal1 ;
  RECT 963.260 1710.800 966.800 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 954.580 1710.800 958.120 1711.920 ;
  LAYER metal4 ;
  RECT 954.580 1710.800 958.120 1711.920 ;
  LAYER metal3 ;
  RECT 954.580 1710.800 958.120 1711.920 ;
  LAYER metal2 ;
  RECT 954.580 1710.800 958.120 1711.920 ;
  LAYER metal1 ;
  RECT 954.580 1710.800 958.120 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 945.900 1710.800 949.440 1711.920 ;
  LAYER metal4 ;
  RECT 945.900 1710.800 949.440 1711.920 ;
  LAYER metal3 ;
  RECT 945.900 1710.800 949.440 1711.920 ;
  LAYER metal2 ;
  RECT 945.900 1710.800 949.440 1711.920 ;
  LAYER metal1 ;
  RECT 945.900 1710.800 949.440 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 937.220 1710.800 940.760 1711.920 ;
  LAYER metal4 ;
  RECT 937.220 1710.800 940.760 1711.920 ;
  LAYER metal3 ;
  RECT 937.220 1710.800 940.760 1711.920 ;
  LAYER metal2 ;
  RECT 937.220 1710.800 940.760 1711.920 ;
  LAYER metal1 ;
  RECT 937.220 1710.800 940.760 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 879.560 1710.800 883.100 1711.920 ;
  LAYER metal4 ;
  RECT 879.560 1710.800 883.100 1711.920 ;
  LAYER metal3 ;
  RECT 879.560 1710.800 883.100 1711.920 ;
  LAYER metal2 ;
  RECT 879.560 1710.800 883.100 1711.920 ;
  LAYER metal1 ;
  RECT 879.560 1710.800 883.100 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 865.300 1710.800 868.840 1711.920 ;
  LAYER metal4 ;
  RECT 865.300 1710.800 868.840 1711.920 ;
  LAYER metal3 ;
  RECT 865.300 1710.800 868.840 1711.920 ;
  LAYER metal2 ;
  RECT 865.300 1710.800 868.840 1711.920 ;
  LAYER metal1 ;
  RECT 865.300 1710.800 868.840 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 856.620 1710.800 860.160 1711.920 ;
  LAYER metal4 ;
  RECT 856.620 1710.800 860.160 1711.920 ;
  LAYER metal3 ;
  RECT 856.620 1710.800 860.160 1711.920 ;
  LAYER metal2 ;
  RECT 856.620 1710.800 860.160 1711.920 ;
  LAYER metal1 ;
  RECT 856.620 1710.800 860.160 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 847.940 1710.800 851.480 1711.920 ;
  LAYER metal4 ;
  RECT 847.940 1710.800 851.480 1711.920 ;
  LAYER metal3 ;
  RECT 847.940 1710.800 851.480 1711.920 ;
  LAYER metal2 ;
  RECT 847.940 1710.800 851.480 1711.920 ;
  LAYER metal1 ;
  RECT 847.940 1710.800 851.480 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 839.260 1710.800 842.800 1711.920 ;
  LAYER metal4 ;
  RECT 839.260 1710.800 842.800 1711.920 ;
  LAYER metal3 ;
  RECT 839.260 1710.800 842.800 1711.920 ;
  LAYER metal2 ;
  RECT 839.260 1710.800 842.800 1711.920 ;
  LAYER metal1 ;
  RECT 839.260 1710.800 842.800 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 830.580 1710.800 834.120 1711.920 ;
  LAYER metal4 ;
  RECT 830.580 1710.800 834.120 1711.920 ;
  LAYER metal3 ;
  RECT 830.580 1710.800 834.120 1711.920 ;
  LAYER metal2 ;
  RECT 830.580 1710.800 834.120 1711.920 ;
  LAYER metal1 ;
  RECT 830.580 1710.800 834.120 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 787.180 1710.800 790.720 1711.920 ;
  LAYER metal4 ;
  RECT 787.180 1710.800 790.720 1711.920 ;
  LAYER metal3 ;
  RECT 787.180 1710.800 790.720 1711.920 ;
  LAYER metal2 ;
  RECT 787.180 1710.800 790.720 1711.920 ;
  LAYER metal1 ;
  RECT 787.180 1710.800 790.720 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 778.500 1710.800 782.040 1711.920 ;
  LAYER metal4 ;
  RECT 778.500 1710.800 782.040 1711.920 ;
  LAYER metal3 ;
  RECT 778.500 1710.800 782.040 1711.920 ;
  LAYER metal2 ;
  RECT 778.500 1710.800 782.040 1711.920 ;
  LAYER metal1 ;
  RECT 778.500 1710.800 782.040 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 769.820 1710.800 773.360 1711.920 ;
  LAYER metal4 ;
  RECT 769.820 1710.800 773.360 1711.920 ;
  LAYER metal3 ;
  RECT 769.820 1710.800 773.360 1711.920 ;
  LAYER metal2 ;
  RECT 769.820 1710.800 773.360 1711.920 ;
  LAYER metal1 ;
  RECT 769.820 1710.800 773.360 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 761.140 1710.800 764.680 1711.920 ;
  LAYER metal4 ;
  RECT 761.140 1710.800 764.680 1711.920 ;
  LAYER metal3 ;
  RECT 761.140 1710.800 764.680 1711.920 ;
  LAYER metal2 ;
  RECT 761.140 1710.800 764.680 1711.920 ;
  LAYER metal1 ;
  RECT 761.140 1710.800 764.680 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 752.460 1710.800 756.000 1711.920 ;
  LAYER metal4 ;
  RECT 752.460 1710.800 756.000 1711.920 ;
  LAYER metal3 ;
  RECT 752.460 1710.800 756.000 1711.920 ;
  LAYER metal2 ;
  RECT 752.460 1710.800 756.000 1711.920 ;
  LAYER metal1 ;
  RECT 752.460 1710.800 756.000 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 743.780 1710.800 747.320 1711.920 ;
  LAYER metal4 ;
  RECT 743.780 1710.800 747.320 1711.920 ;
  LAYER metal3 ;
  RECT 743.780 1710.800 747.320 1711.920 ;
  LAYER metal2 ;
  RECT 743.780 1710.800 747.320 1711.920 ;
  LAYER metal1 ;
  RECT 743.780 1710.800 747.320 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 700.380 1710.800 703.920 1711.920 ;
  LAYER metal4 ;
  RECT 700.380 1710.800 703.920 1711.920 ;
  LAYER metal3 ;
  RECT 700.380 1710.800 703.920 1711.920 ;
  LAYER metal2 ;
  RECT 700.380 1710.800 703.920 1711.920 ;
  LAYER metal1 ;
  RECT 700.380 1710.800 703.920 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 691.700 1710.800 695.240 1711.920 ;
  LAYER metal4 ;
  RECT 691.700 1710.800 695.240 1711.920 ;
  LAYER metal3 ;
  RECT 691.700 1710.800 695.240 1711.920 ;
  LAYER metal2 ;
  RECT 691.700 1710.800 695.240 1711.920 ;
  LAYER metal1 ;
  RECT 691.700 1710.800 695.240 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 683.020 1710.800 686.560 1711.920 ;
  LAYER metal4 ;
  RECT 683.020 1710.800 686.560 1711.920 ;
  LAYER metal3 ;
  RECT 683.020 1710.800 686.560 1711.920 ;
  LAYER metal2 ;
  RECT 683.020 1710.800 686.560 1711.920 ;
  LAYER metal1 ;
  RECT 683.020 1710.800 686.560 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 674.340 1710.800 677.880 1711.920 ;
  LAYER metal4 ;
  RECT 674.340 1710.800 677.880 1711.920 ;
  LAYER metal3 ;
  RECT 674.340 1710.800 677.880 1711.920 ;
  LAYER metal2 ;
  RECT 674.340 1710.800 677.880 1711.920 ;
  LAYER metal1 ;
  RECT 674.340 1710.800 677.880 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 665.660 1710.800 669.200 1711.920 ;
  LAYER metal4 ;
  RECT 665.660 1710.800 669.200 1711.920 ;
  LAYER metal3 ;
  RECT 665.660 1710.800 669.200 1711.920 ;
  LAYER metal2 ;
  RECT 665.660 1710.800 669.200 1711.920 ;
  LAYER metal1 ;
  RECT 665.660 1710.800 669.200 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 656.980 1710.800 660.520 1711.920 ;
  LAYER metal4 ;
  RECT 656.980 1710.800 660.520 1711.920 ;
  LAYER metal3 ;
  RECT 656.980 1710.800 660.520 1711.920 ;
  LAYER metal2 ;
  RECT 656.980 1710.800 660.520 1711.920 ;
  LAYER metal1 ;
  RECT 656.980 1710.800 660.520 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 613.580 1710.800 617.120 1711.920 ;
  LAYER metal4 ;
  RECT 613.580 1710.800 617.120 1711.920 ;
  LAYER metal3 ;
  RECT 613.580 1710.800 617.120 1711.920 ;
  LAYER metal2 ;
  RECT 613.580 1710.800 617.120 1711.920 ;
  LAYER metal1 ;
  RECT 613.580 1710.800 617.120 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 604.900 1710.800 608.440 1711.920 ;
  LAYER metal4 ;
  RECT 604.900 1710.800 608.440 1711.920 ;
  LAYER metal3 ;
  RECT 604.900 1710.800 608.440 1711.920 ;
  LAYER metal2 ;
  RECT 604.900 1710.800 608.440 1711.920 ;
  LAYER metal1 ;
  RECT 604.900 1710.800 608.440 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 596.220 1710.800 599.760 1711.920 ;
  LAYER metal4 ;
  RECT 596.220 1710.800 599.760 1711.920 ;
  LAYER metal3 ;
  RECT 596.220 1710.800 599.760 1711.920 ;
  LAYER metal2 ;
  RECT 596.220 1710.800 599.760 1711.920 ;
  LAYER metal1 ;
  RECT 596.220 1710.800 599.760 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 587.540 1710.800 591.080 1711.920 ;
  LAYER metal4 ;
  RECT 587.540 1710.800 591.080 1711.920 ;
  LAYER metal3 ;
  RECT 587.540 1710.800 591.080 1711.920 ;
  LAYER metal2 ;
  RECT 587.540 1710.800 591.080 1711.920 ;
  LAYER metal1 ;
  RECT 587.540 1710.800 591.080 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 578.860 1710.800 582.400 1711.920 ;
  LAYER metal4 ;
  RECT 578.860 1710.800 582.400 1711.920 ;
  LAYER metal3 ;
  RECT 578.860 1710.800 582.400 1711.920 ;
  LAYER metal2 ;
  RECT 578.860 1710.800 582.400 1711.920 ;
  LAYER metal1 ;
  RECT 578.860 1710.800 582.400 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 570.180 1710.800 573.720 1711.920 ;
  LAYER metal4 ;
  RECT 570.180 1710.800 573.720 1711.920 ;
  LAYER metal3 ;
  RECT 570.180 1710.800 573.720 1711.920 ;
  LAYER metal2 ;
  RECT 570.180 1710.800 573.720 1711.920 ;
  LAYER metal1 ;
  RECT 570.180 1710.800 573.720 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 526.780 1710.800 530.320 1711.920 ;
  LAYER metal4 ;
  RECT 526.780 1710.800 530.320 1711.920 ;
  LAYER metal3 ;
  RECT 526.780 1710.800 530.320 1711.920 ;
  LAYER metal2 ;
  RECT 526.780 1710.800 530.320 1711.920 ;
  LAYER metal1 ;
  RECT 526.780 1710.800 530.320 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 518.100 1710.800 521.640 1711.920 ;
  LAYER metal4 ;
  RECT 518.100 1710.800 521.640 1711.920 ;
  LAYER metal3 ;
  RECT 518.100 1710.800 521.640 1711.920 ;
  LAYER metal2 ;
  RECT 518.100 1710.800 521.640 1711.920 ;
  LAYER metal1 ;
  RECT 518.100 1710.800 521.640 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 509.420 1710.800 512.960 1711.920 ;
  LAYER metal4 ;
  RECT 509.420 1710.800 512.960 1711.920 ;
  LAYER metal3 ;
  RECT 509.420 1710.800 512.960 1711.920 ;
  LAYER metal2 ;
  RECT 509.420 1710.800 512.960 1711.920 ;
  LAYER metal1 ;
  RECT 509.420 1710.800 512.960 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 500.740 1710.800 504.280 1711.920 ;
  LAYER metal4 ;
  RECT 500.740 1710.800 504.280 1711.920 ;
  LAYER metal3 ;
  RECT 500.740 1710.800 504.280 1711.920 ;
  LAYER metal2 ;
  RECT 500.740 1710.800 504.280 1711.920 ;
  LAYER metal1 ;
  RECT 500.740 1710.800 504.280 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 492.060 1710.800 495.600 1711.920 ;
  LAYER metal4 ;
  RECT 492.060 1710.800 495.600 1711.920 ;
  LAYER metal3 ;
  RECT 492.060 1710.800 495.600 1711.920 ;
  LAYER metal2 ;
  RECT 492.060 1710.800 495.600 1711.920 ;
  LAYER metal1 ;
  RECT 492.060 1710.800 495.600 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 478.420 1710.800 481.960 1711.920 ;
  LAYER metal4 ;
  RECT 478.420 1710.800 481.960 1711.920 ;
  LAYER metal3 ;
  RECT 478.420 1710.800 481.960 1711.920 ;
  LAYER metal2 ;
  RECT 478.420 1710.800 481.960 1711.920 ;
  LAYER metal1 ;
  RECT 478.420 1710.800 481.960 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 419.520 1710.800 423.060 1711.920 ;
  LAYER metal4 ;
  RECT 419.520 1710.800 423.060 1711.920 ;
  LAYER metal3 ;
  RECT 419.520 1710.800 423.060 1711.920 ;
  LAYER metal2 ;
  RECT 419.520 1710.800 423.060 1711.920 ;
  LAYER metal1 ;
  RECT 419.520 1710.800 423.060 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 410.840 1710.800 414.380 1711.920 ;
  LAYER metal4 ;
  RECT 410.840 1710.800 414.380 1711.920 ;
  LAYER metal3 ;
  RECT 410.840 1710.800 414.380 1711.920 ;
  LAYER metal2 ;
  RECT 410.840 1710.800 414.380 1711.920 ;
  LAYER metal1 ;
  RECT 410.840 1710.800 414.380 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 402.160 1710.800 405.700 1711.920 ;
  LAYER metal4 ;
  RECT 402.160 1710.800 405.700 1711.920 ;
  LAYER metal3 ;
  RECT 402.160 1710.800 405.700 1711.920 ;
  LAYER metal2 ;
  RECT 402.160 1710.800 405.700 1711.920 ;
  LAYER metal1 ;
  RECT 402.160 1710.800 405.700 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 393.480 1710.800 397.020 1711.920 ;
  LAYER metal4 ;
  RECT 393.480 1710.800 397.020 1711.920 ;
  LAYER metal3 ;
  RECT 393.480 1710.800 397.020 1711.920 ;
  LAYER metal2 ;
  RECT 393.480 1710.800 397.020 1711.920 ;
  LAYER metal1 ;
  RECT 393.480 1710.800 397.020 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 384.800 1710.800 388.340 1711.920 ;
  LAYER metal4 ;
  RECT 384.800 1710.800 388.340 1711.920 ;
  LAYER metal3 ;
  RECT 384.800 1710.800 388.340 1711.920 ;
  LAYER metal2 ;
  RECT 384.800 1710.800 388.340 1711.920 ;
  LAYER metal1 ;
  RECT 384.800 1710.800 388.340 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 376.120 1710.800 379.660 1711.920 ;
  LAYER metal4 ;
  RECT 376.120 1710.800 379.660 1711.920 ;
  LAYER metal3 ;
  RECT 376.120 1710.800 379.660 1711.920 ;
  LAYER metal2 ;
  RECT 376.120 1710.800 379.660 1711.920 ;
  LAYER metal1 ;
  RECT 376.120 1710.800 379.660 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 332.720 1710.800 336.260 1711.920 ;
  LAYER metal4 ;
  RECT 332.720 1710.800 336.260 1711.920 ;
  LAYER metal3 ;
  RECT 332.720 1710.800 336.260 1711.920 ;
  LAYER metal2 ;
  RECT 332.720 1710.800 336.260 1711.920 ;
  LAYER metal1 ;
  RECT 332.720 1710.800 336.260 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 324.040 1710.800 327.580 1711.920 ;
  LAYER metal4 ;
  RECT 324.040 1710.800 327.580 1711.920 ;
  LAYER metal3 ;
  RECT 324.040 1710.800 327.580 1711.920 ;
  LAYER metal2 ;
  RECT 324.040 1710.800 327.580 1711.920 ;
  LAYER metal1 ;
  RECT 324.040 1710.800 327.580 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 315.360 1710.800 318.900 1711.920 ;
  LAYER metal4 ;
  RECT 315.360 1710.800 318.900 1711.920 ;
  LAYER metal3 ;
  RECT 315.360 1710.800 318.900 1711.920 ;
  LAYER metal2 ;
  RECT 315.360 1710.800 318.900 1711.920 ;
  LAYER metal1 ;
  RECT 315.360 1710.800 318.900 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 306.680 1710.800 310.220 1711.920 ;
  LAYER metal4 ;
  RECT 306.680 1710.800 310.220 1711.920 ;
  LAYER metal3 ;
  RECT 306.680 1710.800 310.220 1711.920 ;
  LAYER metal2 ;
  RECT 306.680 1710.800 310.220 1711.920 ;
  LAYER metal1 ;
  RECT 306.680 1710.800 310.220 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 298.000 1710.800 301.540 1711.920 ;
  LAYER metal4 ;
  RECT 298.000 1710.800 301.540 1711.920 ;
  LAYER metal3 ;
  RECT 298.000 1710.800 301.540 1711.920 ;
  LAYER metal2 ;
  RECT 298.000 1710.800 301.540 1711.920 ;
  LAYER metal1 ;
  RECT 298.000 1710.800 301.540 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 289.320 1710.800 292.860 1711.920 ;
  LAYER metal4 ;
  RECT 289.320 1710.800 292.860 1711.920 ;
  LAYER metal3 ;
  RECT 289.320 1710.800 292.860 1711.920 ;
  LAYER metal2 ;
  RECT 289.320 1710.800 292.860 1711.920 ;
  LAYER metal1 ;
  RECT 289.320 1710.800 292.860 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 245.920 1710.800 249.460 1711.920 ;
  LAYER metal4 ;
  RECT 245.920 1710.800 249.460 1711.920 ;
  LAYER metal3 ;
  RECT 245.920 1710.800 249.460 1711.920 ;
  LAYER metal2 ;
  RECT 245.920 1710.800 249.460 1711.920 ;
  LAYER metal1 ;
  RECT 245.920 1710.800 249.460 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 237.240 1710.800 240.780 1711.920 ;
  LAYER metal4 ;
  RECT 237.240 1710.800 240.780 1711.920 ;
  LAYER metal3 ;
  RECT 237.240 1710.800 240.780 1711.920 ;
  LAYER metal2 ;
  RECT 237.240 1710.800 240.780 1711.920 ;
  LAYER metal1 ;
  RECT 237.240 1710.800 240.780 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 228.560 1710.800 232.100 1711.920 ;
  LAYER metal4 ;
  RECT 228.560 1710.800 232.100 1711.920 ;
  LAYER metal3 ;
  RECT 228.560 1710.800 232.100 1711.920 ;
  LAYER metal2 ;
  RECT 228.560 1710.800 232.100 1711.920 ;
  LAYER metal1 ;
  RECT 228.560 1710.800 232.100 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 219.880 1710.800 223.420 1711.920 ;
  LAYER metal4 ;
  RECT 219.880 1710.800 223.420 1711.920 ;
  LAYER metal3 ;
  RECT 219.880 1710.800 223.420 1711.920 ;
  LAYER metal2 ;
  RECT 219.880 1710.800 223.420 1711.920 ;
  LAYER metal1 ;
  RECT 219.880 1710.800 223.420 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 211.200 1710.800 214.740 1711.920 ;
  LAYER metal4 ;
  RECT 211.200 1710.800 214.740 1711.920 ;
  LAYER metal3 ;
  RECT 211.200 1710.800 214.740 1711.920 ;
  LAYER metal2 ;
  RECT 211.200 1710.800 214.740 1711.920 ;
  LAYER metal1 ;
  RECT 211.200 1710.800 214.740 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 202.520 1710.800 206.060 1711.920 ;
  LAYER metal4 ;
  RECT 202.520 1710.800 206.060 1711.920 ;
  LAYER metal3 ;
  RECT 202.520 1710.800 206.060 1711.920 ;
  LAYER metal2 ;
  RECT 202.520 1710.800 206.060 1711.920 ;
  LAYER metal1 ;
  RECT 202.520 1710.800 206.060 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 159.120 1710.800 162.660 1711.920 ;
  LAYER metal4 ;
  RECT 159.120 1710.800 162.660 1711.920 ;
  LAYER metal3 ;
  RECT 159.120 1710.800 162.660 1711.920 ;
  LAYER metal2 ;
  RECT 159.120 1710.800 162.660 1711.920 ;
  LAYER metal1 ;
  RECT 159.120 1710.800 162.660 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 150.440 1710.800 153.980 1711.920 ;
  LAYER metal4 ;
  RECT 150.440 1710.800 153.980 1711.920 ;
  LAYER metal3 ;
  RECT 150.440 1710.800 153.980 1711.920 ;
  LAYER metal2 ;
  RECT 150.440 1710.800 153.980 1711.920 ;
  LAYER metal1 ;
  RECT 150.440 1710.800 153.980 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 141.760 1710.800 145.300 1711.920 ;
  LAYER metal4 ;
  RECT 141.760 1710.800 145.300 1711.920 ;
  LAYER metal3 ;
  RECT 141.760 1710.800 145.300 1711.920 ;
  LAYER metal2 ;
  RECT 141.760 1710.800 145.300 1711.920 ;
  LAYER metal1 ;
  RECT 141.760 1710.800 145.300 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 133.080 1710.800 136.620 1711.920 ;
  LAYER metal4 ;
  RECT 133.080 1710.800 136.620 1711.920 ;
  LAYER metal3 ;
  RECT 133.080 1710.800 136.620 1711.920 ;
  LAYER metal2 ;
  RECT 133.080 1710.800 136.620 1711.920 ;
  LAYER metal1 ;
  RECT 133.080 1710.800 136.620 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 124.400 1710.800 127.940 1711.920 ;
  LAYER metal4 ;
  RECT 124.400 1710.800 127.940 1711.920 ;
  LAYER metal3 ;
  RECT 124.400 1710.800 127.940 1711.920 ;
  LAYER metal2 ;
  RECT 124.400 1710.800 127.940 1711.920 ;
  LAYER metal1 ;
  RECT 124.400 1710.800 127.940 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 115.720 1710.800 119.260 1711.920 ;
  LAYER metal4 ;
  RECT 115.720 1710.800 119.260 1711.920 ;
  LAYER metal3 ;
  RECT 115.720 1710.800 119.260 1711.920 ;
  LAYER metal2 ;
  RECT 115.720 1710.800 119.260 1711.920 ;
  LAYER metal1 ;
  RECT 115.720 1710.800 119.260 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 72.320 1710.800 75.860 1711.920 ;
  LAYER metal4 ;
  RECT 72.320 1710.800 75.860 1711.920 ;
  LAYER metal3 ;
  RECT 72.320 1710.800 75.860 1711.920 ;
  LAYER metal2 ;
  RECT 72.320 1710.800 75.860 1711.920 ;
  LAYER metal1 ;
  RECT 72.320 1710.800 75.860 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 63.640 1710.800 67.180 1711.920 ;
  LAYER metal4 ;
  RECT 63.640 1710.800 67.180 1711.920 ;
  LAYER metal3 ;
  RECT 63.640 1710.800 67.180 1711.920 ;
  LAYER metal2 ;
  RECT 63.640 1710.800 67.180 1711.920 ;
  LAYER metal1 ;
  RECT 63.640 1710.800 67.180 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 54.960 1710.800 58.500 1711.920 ;
  LAYER metal4 ;
  RECT 54.960 1710.800 58.500 1711.920 ;
  LAYER metal3 ;
  RECT 54.960 1710.800 58.500 1711.920 ;
  LAYER metal2 ;
  RECT 54.960 1710.800 58.500 1711.920 ;
  LAYER metal1 ;
  RECT 54.960 1710.800 58.500 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 41.940 1710.800 45.480 1711.920 ;
  LAYER metal4 ;
  RECT 41.940 1710.800 45.480 1711.920 ;
  LAYER metal3 ;
  RECT 41.940 1710.800 45.480 1711.920 ;
  LAYER metal2 ;
  RECT 41.940 1710.800 45.480 1711.920 ;
  LAYER metal1 ;
  RECT 41.940 1710.800 45.480 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 28.300 1710.800 31.840 1711.920 ;
  LAYER metal4 ;
  RECT 28.300 1710.800 31.840 1711.920 ;
  LAYER metal3 ;
  RECT 28.300 1710.800 31.840 1711.920 ;
  LAYER metal2 ;
  RECT 28.300 1710.800 31.840 1711.920 ;
  LAYER metal1 ;
  RECT 28.300 1710.800 31.840 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 14.660 1710.800 18.200 1711.920 ;
  LAYER metal4 ;
  RECT 14.660 1710.800 18.200 1711.920 ;
  LAYER metal3 ;
  RECT 14.660 1710.800 18.200 1711.920 ;
  LAYER metal2 ;
  RECT 14.660 1710.800 18.200 1711.920 ;
  LAYER metal1 ;
  RECT 14.660 1710.800 18.200 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3592.060 0.000 3595.600 1.120 ;
  LAYER metal4 ;
  RECT 3592.060 0.000 3595.600 1.120 ;
  LAYER metal3 ;
  RECT 3592.060 0.000 3595.600 1.120 ;
  LAYER metal2 ;
  RECT 3592.060 0.000 3595.600 1.120 ;
  LAYER metal1 ;
  RECT 3592.060 0.000 3595.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3583.380 0.000 3586.920 1.120 ;
  LAYER metal4 ;
  RECT 3583.380 0.000 3586.920 1.120 ;
  LAYER metal3 ;
  RECT 3583.380 0.000 3586.920 1.120 ;
  LAYER metal2 ;
  RECT 3583.380 0.000 3586.920 1.120 ;
  LAYER metal1 ;
  RECT 3583.380 0.000 3586.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3574.700 0.000 3578.240 1.120 ;
  LAYER metal4 ;
  RECT 3574.700 0.000 3578.240 1.120 ;
  LAYER metal3 ;
  RECT 3574.700 0.000 3578.240 1.120 ;
  LAYER metal2 ;
  RECT 3574.700 0.000 3578.240 1.120 ;
  LAYER metal1 ;
  RECT 3574.700 0.000 3578.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3566.020 0.000 3569.560 1.120 ;
  LAYER metal4 ;
  RECT 3566.020 0.000 3569.560 1.120 ;
  LAYER metal3 ;
  RECT 3566.020 0.000 3569.560 1.120 ;
  LAYER metal2 ;
  RECT 3566.020 0.000 3569.560 1.120 ;
  LAYER metal1 ;
  RECT 3566.020 0.000 3569.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3557.340 0.000 3560.880 1.120 ;
  LAYER metal4 ;
  RECT 3557.340 0.000 3560.880 1.120 ;
  LAYER metal3 ;
  RECT 3557.340 0.000 3560.880 1.120 ;
  LAYER metal2 ;
  RECT 3557.340 0.000 3560.880 1.120 ;
  LAYER metal1 ;
  RECT 3557.340 0.000 3560.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3548.660 0.000 3552.200 1.120 ;
  LAYER metal4 ;
  RECT 3548.660 0.000 3552.200 1.120 ;
  LAYER metal3 ;
  RECT 3548.660 0.000 3552.200 1.120 ;
  LAYER metal2 ;
  RECT 3548.660 0.000 3552.200 1.120 ;
  LAYER metal1 ;
  RECT 3548.660 0.000 3552.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3505.260 0.000 3508.800 1.120 ;
  LAYER metal4 ;
  RECT 3505.260 0.000 3508.800 1.120 ;
  LAYER metal3 ;
  RECT 3505.260 0.000 3508.800 1.120 ;
  LAYER metal2 ;
  RECT 3505.260 0.000 3508.800 1.120 ;
  LAYER metal1 ;
  RECT 3505.260 0.000 3508.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3496.580 0.000 3500.120 1.120 ;
  LAYER metal4 ;
  RECT 3496.580 0.000 3500.120 1.120 ;
  LAYER metal3 ;
  RECT 3496.580 0.000 3500.120 1.120 ;
  LAYER metal2 ;
  RECT 3496.580 0.000 3500.120 1.120 ;
  LAYER metal1 ;
  RECT 3496.580 0.000 3500.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3487.900 0.000 3491.440 1.120 ;
  LAYER metal4 ;
  RECT 3487.900 0.000 3491.440 1.120 ;
  LAYER metal3 ;
  RECT 3487.900 0.000 3491.440 1.120 ;
  LAYER metal2 ;
  RECT 3487.900 0.000 3491.440 1.120 ;
  LAYER metal1 ;
  RECT 3487.900 0.000 3491.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3479.220 0.000 3482.760 1.120 ;
  LAYER metal4 ;
  RECT 3479.220 0.000 3482.760 1.120 ;
  LAYER metal3 ;
  RECT 3479.220 0.000 3482.760 1.120 ;
  LAYER metal2 ;
  RECT 3479.220 0.000 3482.760 1.120 ;
  LAYER metal1 ;
  RECT 3479.220 0.000 3482.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3470.540 0.000 3474.080 1.120 ;
  LAYER metal4 ;
  RECT 3470.540 0.000 3474.080 1.120 ;
  LAYER metal3 ;
  RECT 3470.540 0.000 3474.080 1.120 ;
  LAYER metal2 ;
  RECT 3470.540 0.000 3474.080 1.120 ;
  LAYER metal1 ;
  RECT 3470.540 0.000 3474.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3461.860 0.000 3465.400 1.120 ;
  LAYER metal4 ;
  RECT 3461.860 0.000 3465.400 1.120 ;
  LAYER metal3 ;
  RECT 3461.860 0.000 3465.400 1.120 ;
  LAYER metal2 ;
  RECT 3461.860 0.000 3465.400 1.120 ;
  LAYER metal1 ;
  RECT 3461.860 0.000 3465.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3418.460 0.000 3422.000 1.120 ;
  LAYER metal4 ;
  RECT 3418.460 0.000 3422.000 1.120 ;
  LAYER metal3 ;
  RECT 3418.460 0.000 3422.000 1.120 ;
  LAYER metal2 ;
  RECT 3418.460 0.000 3422.000 1.120 ;
  LAYER metal1 ;
  RECT 3418.460 0.000 3422.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3409.780 0.000 3413.320 1.120 ;
  LAYER metal4 ;
  RECT 3409.780 0.000 3413.320 1.120 ;
  LAYER metal3 ;
  RECT 3409.780 0.000 3413.320 1.120 ;
  LAYER metal2 ;
  RECT 3409.780 0.000 3413.320 1.120 ;
  LAYER metal1 ;
  RECT 3409.780 0.000 3413.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3401.100 0.000 3404.640 1.120 ;
  LAYER metal4 ;
  RECT 3401.100 0.000 3404.640 1.120 ;
  LAYER metal3 ;
  RECT 3401.100 0.000 3404.640 1.120 ;
  LAYER metal2 ;
  RECT 3401.100 0.000 3404.640 1.120 ;
  LAYER metal1 ;
  RECT 3401.100 0.000 3404.640 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3392.420 0.000 3395.960 1.120 ;
  LAYER metal4 ;
  RECT 3392.420 0.000 3395.960 1.120 ;
  LAYER metal3 ;
  RECT 3392.420 0.000 3395.960 1.120 ;
  LAYER metal2 ;
  RECT 3392.420 0.000 3395.960 1.120 ;
  LAYER metal1 ;
  RECT 3392.420 0.000 3395.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3383.740 0.000 3387.280 1.120 ;
  LAYER metal4 ;
  RECT 3383.740 0.000 3387.280 1.120 ;
  LAYER metal3 ;
  RECT 3383.740 0.000 3387.280 1.120 ;
  LAYER metal2 ;
  RECT 3383.740 0.000 3387.280 1.120 ;
  LAYER metal1 ;
  RECT 3383.740 0.000 3387.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3375.060 0.000 3378.600 1.120 ;
  LAYER metal4 ;
  RECT 3375.060 0.000 3378.600 1.120 ;
  LAYER metal3 ;
  RECT 3375.060 0.000 3378.600 1.120 ;
  LAYER metal2 ;
  RECT 3375.060 0.000 3378.600 1.120 ;
  LAYER metal1 ;
  RECT 3375.060 0.000 3378.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3331.660 0.000 3335.200 1.120 ;
  LAYER metal4 ;
  RECT 3331.660 0.000 3335.200 1.120 ;
  LAYER metal3 ;
  RECT 3331.660 0.000 3335.200 1.120 ;
  LAYER metal2 ;
  RECT 3331.660 0.000 3335.200 1.120 ;
  LAYER metal1 ;
  RECT 3331.660 0.000 3335.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3322.980 0.000 3326.520 1.120 ;
  LAYER metal4 ;
  RECT 3322.980 0.000 3326.520 1.120 ;
  LAYER metal3 ;
  RECT 3322.980 0.000 3326.520 1.120 ;
  LAYER metal2 ;
  RECT 3322.980 0.000 3326.520 1.120 ;
  LAYER metal1 ;
  RECT 3322.980 0.000 3326.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3314.300 0.000 3317.840 1.120 ;
  LAYER metal4 ;
  RECT 3314.300 0.000 3317.840 1.120 ;
  LAYER metal3 ;
  RECT 3314.300 0.000 3317.840 1.120 ;
  LAYER metal2 ;
  RECT 3314.300 0.000 3317.840 1.120 ;
  LAYER metal1 ;
  RECT 3314.300 0.000 3317.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3305.620 0.000 3309.160 1.120 ;
  LAYER metal4 ;
  RECT 3305.620 0.000 3309.160 1.120 ;
  LAYER metal3 ;
  RECT 3305.620 0.000 3309.160 1.120 ;
  LAYER metal2 ;
  RECT 3305.620 0.000 3309.160 1.120 ;
  LAYER metal1 ;
  RECT 3305.620 0.000 3309.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3296.940 0.000 3300.480 1.120 ;
  LAYER metal4 ;
  RECT 3296.940 0.000 3300.480 1.120 ;
  LAYER metal3 ;
  RECT 3296.940 0.000 3300.480 1.120 ;
  LAYER metal2 ;
  RECT 3296.940 0.000 3300.480 1.120 ;
  LAYER metal1 ;
  RECT 3296.940 0.000 3300.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3288.260 0.000 3291.800 1.120 ;
  LAYER metal4 ;
  RECT 3288.260 0.000 3291.800 1.120 ;
  LAYER metal3 ;
  RECT 3288.260 0.000 3291.800 1.120 ;
  LAYER metal2 ;
  RECT 3288.260 0.000 3291.800 1.120 ;
  LAYER metal1 ;
  RECT 3288.260 0.000 3291.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3244.860 0.000 3248.400 1.120 ;
  LAYER metal4 ;
  RECT 3244.860 0.000 3248.400 1.120 ;
  LAYER metal3 ;
  RECT 3244.860 0.000 3248.400 1.120 ;
  LAYER metal2 ;
  RECT 3244.860 0.000 3248.400 1.120 ;
  LAYER metal1 ;
  RECT 3244.860 0.000 3248.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3236.180 0.000 3239.720 1.120 ;
  LAYER metal4 ;
  RECT 3236.180 0.000 3239.720 1.120 ;
  LAYER metal3 ;
  RECT 3236.180 0.000 3239.720 1.120 ;
  LAYER metal2 ;
  RECT 3236.180 0.000 3239.720 1.120 ;
  LAYER metal1 ;
  RECT 3236.180 0.000 3239.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3227.500 0.000 3231.040 1.120 ;
  LAYER metal4 ;
  RECT 3227.500 0.000 3231.040 1.120 ;
  LAYER metal3 ;
  RECT 3227.500 0.000 3231.040 1.120 ;
  LAYER metal2 ;
  RECT 3227.500 0.000 3231.040 1.120 ;
  LAYER metal1 ;
  RECT 3227.500 0.000 3231.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3218.820 0.000 3222.360 1.120 ;
  LAYER metal4 ;
  RECT 3218.820 0.000 3222.360 1.120 ;
  LAYER metal3 ;
  RECT 3218.820 0.000 3222.360 1.120 ;
  LAYER metal2 ;
  RECT 3218.820 0.000 3222.360 1.120 ;
  LAYER metal1 ;
  RECT 3218.820 0.000 3222.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3205.800 0.000 3209.340 1.120 ;
  LAYER metal4 ;
  RECT 3205.800 0.000 3209.340 1.120 ;
  LAYER metal3 ;
  RECT 3205.800 0.000 3209.340 1.120 ;
  LAYER metal2 ;
  RECT 3205.800 0.000 3209.340 1.120 ;
  LAYER metal1 ;
  RECT 3205.800 0.000 3209.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3192.160 0.000 3195.700 1.120 ;
  LAYER metal4 ;
  RECT 3192.160 0.000 3195.700 1.120 ;
  LAYER metal3 ;
  RECT 3192.160 0.000 3195.700 1.120 ;
  LAYER metal2 ;
  RECT 3192.160 0.000 3195.700 1.120 ;
  LAYER metal1 ;
  RECT 3192.160 0.000 3195.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3138.220 0.000 3141.760 1.120 ;
  LAYER metal4 ;
  RECT 3138.220 0.000 3141.760 1.120 ;
  LAYER metal3 ;
  RECT 3138.220 0.000 3141.760 1.120 ;
  LAYER metal2 ;
  RECT 3138.220 0.000 3141.760 1.120 ;
  LAYER metal1 ;
  RECT 3138.220 0.000 3141.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3129.540 0.000 3133.080 1.120 ;
  LAYER metal4 ;
  RECT 3129.540 0.000 3133.080 1.120 ;
  LAYER metal3 ;
  RECT 3129.540 0.000 3133.080 1.120 ;
  LAYER metal2 ;
  RECT 3129.540 0.000 3133.080 1.120 ;
  LAYER metal1 ;
  RECT 3129.540 0.000 3133.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3120.860 0.000 3124.400 1.120 ;
  LAYER metal4 ;
  RECT 3120.860 0.000 3124.400 1.120 ;
  LAYER metal3 ;
  RECT 3120.860 0.000 3124.400 1.120 ;
  LAYER metal2 ;
  RECT 3120.860 0.000 3124.400 1.120 ;
  LAYER metal1 ;
  RECT 3120.860 0.000 3124.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3112.180 0.000 3115.720 1.120 ;
  LAYER metal4 ;
  RECT 3112.180 0.000 3115.720 1.120 ;
  LAYER metal3 ;
  RECT 3112.180 0.000 3115.720 1.120 ;
  LAYER metal2 ;
  RECT 3112.180 0.000 3115.720 1.120 ;
  LAYER metal1 ;
  RECT 3112.180 0.000 3115.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3103.500 0.000 3107.040 1.120 ;
  LAYER metal4 ;
  RECT 3103.500 0.000 3107.040 1.120 ;
  LAYER metal3 ;
  RECT 3103.500 0.000 3107.040 1.120 ;
  LAYER metal2 ;
  RECT 3103.500 0.000 3107.040 1.120 ;
  LAYER metal1 ;
  RECT 3103.500 0.000 3107.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3094.820 0.000 3098.360 1.120 ;
  LAYER metal4 ;
  RECT 3094.820 0.000 3098.360 1.120 ;
  LAYER metal3 ;
  RECT 3094.820 0.000 3098.360 1.120 ;
  LAYER metal2 ;
  RECT 3094.820 0.000 3098.360 1.120 ;
  LAYER metal1 ;
  RECT 3094.820 0.000 3098.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3051.420 0.000 3054.960 1.120 ;
  LAYER metal4 ;
  RECT 3051.420 0.000 3054.960 1.120 ;
  LAYER metal3 ;
  RECT 3051.420 0.000 3054.960 1.120 ;
  LAYER metal2 ;
  RECT 3051.420 0.000 3054.960 1.120 ;
  LAYER metal1 ;
  RECT 3051.420 0.000 3054.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3042.740 0.000 3046.280 1.120 ;
  LAYER metal4 ;
  RECT 3042.740 0.000 3046.280 1.120 ;
  LAYER metal3 ;
  RECT 3042.740 0.000 3046.280 1.120 ;
  LAYER metal2 ;
  RECT 3042.740 0.000 3046.280 1.120 ;
  LAYER metal1 ;
  RECT 3042.740 0.000 3046.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3034.060 0.000 3037.600 1.120 ;
  LAYER metal4 ;
  RECT 3034.060 0.000 3037.600 1.120 ;
  LAYER metal3 ;
  RECT 3034.060 0.000 3037.600 1.120 ;
  LAYER metal2 ;
  RECT 3034.060 0.000 3037.600 1.120 ;
  LAYER metal1 ;
  RECT 3034.060 0.000 3037.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3025.380 0.000 3028.920 1.120 ;
  LAYER metal4 ;
  RECT 3025.380 0.000 3028.920 1.120 ;
  LAYER metal3 ;
  RECT 3025.380 0.000 3028.920 1.120 ;
  LAYER metal2 ;
  RECT 3025.380 0.000 3028.920 1.120 ;
  LAYER metal1 ;
  RECT 3025.380 0.000 3028.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3016.700 0.000 3020.240 1.120 ;
  LAYER metal4 ;
  RECT 3016.700 0.000 3020.240 1.120 ;
  LAYER metal3 ;
  RECT 3016.700 0.000 3020.240 1.120 ;
  LAYER metal2 ;
  RECT 3016.700 0.000 3020.240 1.120 ;
  LAYER metal1 ;
  RECT 3016.700 0.000 3020.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3008.020 0.000 3011.560 1.120 ;
  LAYER metal4 ;
  RECT 3008.020 0.000 3011.560 1.120 ;
  LAYER metal3 ;
  RECT 3008.020 0.000 3011.560 1.120 ;
  LAYER metal2 ;
  RECT 3008.020 0.000 3011.560 1.120 ;
  LAYER metal1 ;
  RECT 3008.020 0.000 3011.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2964.620 0.000 2968.160 1.120 ;
  LAYER metal4 ;
  RECT 2964.620 0.000 2968.160 1.120 ;
  LAYER metal3 ;
  RECT 2964.620 0.000 2968.160 1.120 ;
  LAYER metal2 ;
  RECT 2964.620 0.000 2968.160 1.120 ;
  LAYER metal1 ;
  RECT 2964.620 0.000 2968.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2955.940 0.000 2959.480 1.120 ;
  LAYER metal4 ;
  RECT 2955.940 0.000 2959.480 1.120 ;
  LAYER metal3 ;
  RECT 2955.940 0.000 2959.480 1.120 ;
  LAYER metal2 ;
  RECT 2955.940 0.000 2959.480 1.120 ;
  LAYER metal1 ;
  RECT 2955.940 0.000 2959.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2947.260 0.000 2950.800 1.120 ;
  LAYER metal4 ;
  RECT 2947.260 0.000 2950.800 1.120 ;
  LAYER metal3 ;
  RECT 2947.260 0.000 2950.800 1.120 ;
  LAYER metal2 ;
  RECT 2947.260 0.000 2950.800 1.120 ;
  LAYER metal1 ;
  RECT 2947.260 0.000 2950.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2938.580 0.000 2942.120 1.120 ;
  LAYER metal4 ;
  RECT 2938.580 0.000 2942.120 1.120 ;
  LAYER metal3 ;
  RECT 2938.580 0.000 2942.120 1.120 ;
  LAYER metal2 ;
  RECT 2938.580 0.000 2942.120 1.120 ;
  LAYER metal1 ;
  RECT 2938.580 0.000 2942.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2929.900 0.000 2933.440 1.120 ;
  LAYER metal4 ;
  RECT 2929.900 0.000 2933.440 1.120 ;
  LAYER metal3 ;
  RECT 2929.900 0.000 2933.440 1.120 ;
  LAYER metal2 ;
  RECT 2929.900 0.000 2933.440 1.120 ;
  LAYER metal1 ;
  RECT 2929.900 0.000 2933.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2921.220 0.000 2924.760 1.120 ;
  LAYER metal4 ;
  RECT 2921.220 0.000 2924.760 1.120 ;
  LAYER metal3 ;
  RECT 2921.220 0.000 2924.760 1.120 ;
  LAYER metal2 ;
  RECT 2921.220 0.000 2924.760 1.120 ;
  LAYER metal1 ;
  RECT 2921.220 0.000 2924.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2877.820 0.000 2881.360 1.120 ;
  LAYER metal4 ;
  RECT 2877.820 0.000 2881.360 1.120 ;
  LAYER metal3 ;
  RECT 2877.820 0.000 2881.360 1.120 ;
  LAYER metal2 ;
  RECT 2877.820 0.000 2881.360 1.120 ;
  LAYER metal1 ;
  RECT 2877.820 0.000 2881.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2869.140 0.000 2872.680 1.120 ;
  LAYER metal4 ;
  RECT 2869.140 0.000 2872.680 1.120 ;
  LAYER metal3 ;
  RECT 2869.140 0.000 2872.680 1.120 ;
  LAYER metal2 ;
  RECT 2869.140 0.000 2872.680 1.120 ;
  LAYER metal1 ;
  RECT 2869.140 0.000 2872.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2860.460 0.000 2864.000 1.120 ;
  LAYER metal4 ;
  RECT 2860.460 0.000 2864.000 1.120 ;
  LAYER metal3 ;
  RECT 2860.460 0.000 2864.000 1.120 ;
  LAYER metal2 ;
  RECT 2860.460 0.000 2864.000 1.120 ;
  LAYER metal1 ;
  RECT 2860.460 0.000 2864.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2851.780 0.000 2855.320 1.120 ;
  LAYER metal4 ;
  RECT 2851.780 0.000 2855.320 1.120 ;
  LAYER metal3 ;
  RECT 2851.780 0.000 2855.320 1.120 ;
  LAYER metal2 ;
  RECT 2851.780 0.000 2855.320 1.120 ;
  LAYER metal1 ;
  RECT 2851.780 0.000 2855.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2843.100 0.000 2846.640 1.120 ;
  LAYER metal4 ;
  RECT 2843.100 0.000 2846.640 1.120 ;
  LAYER metal3 ;
  RECT 2843.100 0.000 2846.640 1.120 ;
  LAYER metal2 ;
  RECT 2843.100 0.000 2846.640 1.120 ;
  LAYER metal1 ;
  RECT 2843.100 0.000 2846.640 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2834.420 0.000 2837.960 1.120 ;
  LAYER metal4 ;
  RECT 2834.420 0.000 2837.960 1.120 ;
  LAYER metal3 ;
  RECT 2834.420 0.000 2837.960 1.120 ;
  LAYER metal2 ;
  RECT 2834.420 0.000 2837.960 1.120 ;
  LAYER metal1 ;
  RECT 2834.420 0.000 2837.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2791.020 0.000 2794.560 1.120 ;
  LAYER metal4 ;
  RECT 2791.020 0.000 2794.560 1.120 ;
  LAYER metal3 ;
  RECT 2791.020 0.000 2794.560 1.120 ;
  LAYER metal2 ;
  RECT 2791.020 0.000 2794.560 1.120 ;
  LAYER metal1 ;
  RECT 2791.020 0.000 2794.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2782.340 0.000 2785.880 1.120 ;
  LAYER metal4 ;
  RECT 2782.340 0.000 2785.880 1.120 ;
  LAYER metal3 ;
  RECT 2782.340 0.000 2785.880 1.120 ;
  LAYER metal2 ;
  RECT 2782.340 0.000 2785.880 1.120 ;
  LAYER metal1 ;
  RECT 2782.340 0.000 2785.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2769.320 0.000 2772.860 1.120 ;
  LAYER metal4 ;
  RECT 2769.320 0.000 2772.860 1.120 ;
  LAYER metal3 ;
  RECT 2769.320 0.000 2772.860 1.120 ;
  LAYER metal2 ;
  RECT 2769.320 0.000 2772.860 1.120 ;
  LAYER metal1 ;
  RECT 2769.320 0.000 2772.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2755.680 0.000 2759.220 1.120 ;
  LAYER metal4 ;
  RECT 2755.680 0.000 2759.220 1.120 ;
  LAYER metal3 ;
  RECT 2755.680 0.000 2759.220 1.120 ;
  LAYER metal2 ;
  RECT 2755.680 0.000 2759.220 1.120 ;
  LAYER metal1 ;
  RECT 2755.680 0.000 2759.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2742.040 0.000 2745.580 1.120 ;
  LAYER metal4 ;
  RECT 2742.040 0.000 2745.580 1.120 ;
  LAYER metal3 ;
  RECT 2742.040 0.000 2745.580 1.120 ;
  LAYER metal2 ;
  RECT 2742.040 0.000 2745.580 1.120 ;
  LAYER metal1 ;
  RECT 2742.040 0.000 2745.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2727.780 0.000 2731.320 1.120 ;
  LAYER metal4 ;
  RECT 2727.780 0.000 2731.320 1.120 ;
  LAYER metal3 ;
  RECT 2727.780 0.000 2731.320 1.120 ;
  LAYER metal2 ;
  RECT 2727.780 0.000 2731.320 1.120 ;
  LAYER metal1 ;
  RECT 2727.780 0.000 2731.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2684.380 0.000 2687.920 1.120 ;
  LAYER metal4 ;
  RECT 2684.380 0.000 2687.920 1.120 ;
  LAYER metal3 ;
  RECT 2684.380 0.000 2687.920 1.120 ;
  LAYER metal2 ;
  RECT 2684.380 0.000 2687.920 1.120 ;
  LAYER metal1 ;
  RECT 2684.380 0.000 2687.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2675.700 0.000 2679.240 1.120 ;
  LAYER metal4 ;
  RECT 2675.700 0.000 2679.240 1.120 ;
  LAYER metal3 ;
  RECT 2675.700 0.000 2679.240 1.120 ;
  LAYER metal2 ;
  RECT 2675.700 0.000 2679.240 1.120 ;
  LAYER metal1 ;
  RECT 2675.700 0.000 2679.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2667.020 0.000 2670.560 1.120 ;
  LAYER metal4 ;
  RECT 2667.020 0.000 2670.560 1.120 ;
  LAYER metal3 ;
  RECT 2667.020 0.000 2670.560 1.120 ;
  LAYER metal2 ;
  RECT 2667.020 0.000 2670.560 1.120 ;
  LAYER metal1 ;
  RECT 2667.020 0.000 2670.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2658.340 0.000 2661.880 1.120 ;
  LAYER metal4 ;
  RECT 2658.340 0.000 2661.880 1.120 ;
  LAYER metal3 ;
  RECT 2658.340 0.000 2661.880 1.120 ;
  LAYER metal2 ;
  RECT 2658.340 0.000 2661.880 1.120 ;
  LAYER metal1 ;
  RECT 2658.340 0.000 2661.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2649.660 0.000 2653.200 1.120 ;
  LAYER metal4 ;
  RECT 2649.660 0.000 2653.200 1.120 ;
  LAYER metal3 ;
  RECT 2649.660 0.000 2653.200 1.120 ;
  LAYER metal2 ;
  RECT 2649.660 0.000 2653.200 1.120 ;
  LAYER metal1 ;
  RECT 2649.660 0.000 2653.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2640.980 0.000 2644.520 1.120 ;
  LAYER metal4 ;
  RECT 2640.980 0.000 2644.520 1.120 ;
  LAYER metal3 ;
  RECT 2640.980 0.000 2644.520 1.120 ;
  LAYER metal2 ;
  RECT 2640.980 0.000 2644.520 1.120 ;
  LAYER metal1 ;
  RECT 2640.980 0.000 2644.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2597.580 0.000 2601.120 1.120 ;
  LAYER metal4 ;
  RECT 2597.580 0.000 2601.120 1.120 ;
  LAYER metal3 ;
  RECT 2597.580 0.000 2601.120 1.120 ;
  LAYER metal2 ;
  RECT 2597.580 0.000 2601.120 1.120 ;
  LAYER metal1 ;
  RECT 2597.580 0.000 2601.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2588.900 0.000 2592.440 1.120 ;
  LAYER metal4 ;
  RECT 2588.900 0.000 2592.440 1.120 ;
  LAYER metal3 ;
  RECT 2588.900 0.000 2592.440 1.120 ;
  LAYER metal2 ;
  RECT 2588.900 0.000 2592.440 1.120 ;
  LAYER metal1 ;
  RECT 2588.900 0.000 2592.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2580.220 0.000 2583.760 1.120 ;
  LAYER metal4 ;
  RECT 2580.220 0.000 2583.760 1.120 ;
  LAYER metal3 ;
  RECT 2580.220 0.000 2583.760 1.120 ;
  LAYER metal2 ;
  RECT 2580.220 0.000 2583.760 1.120 ;
  LAYER metal1 ;
  RECT 2580.220 0.000 2583.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2571.540 0.000 2575.080 1.120 ;
  LAYER metal4 ;
  RECT 2571.540 0.000 2575.080 1.120 ;
  LAYER metal3 ;
  RECT 2571.540 0.000 2575.080 1.120 ;
  LAYER metal2 ;
  RECT 2571.540 0.000 2575.080 1.120 ;
  LAYER metal1 ;
  RECT 2571.540 0.000 2575.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2562.860 0.000 2566.400 1.120 ;
  LAYER metal4 ;
  RECT 2562.860 0.000 2566.400 1.120 ;
  LAYER metal3 ;
  RECT 2562.860 0.000 2566.400 1.120 ;
  LAYER metal2 ;
  RECT 2562.860 0.000 2566.400 1.120 ;
  LAYER metal1 ;
  RECT 2562.860 0.000 2566.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2554.180 0.000 2557.720 1.120 ;
  LAYER metal4 ;
  RECT 2554.180 0.000 2557.720 1.120 ;
  LAYER metal3 ;
  RECT 2554.180 0.000 2557.720 1.120 ;
  LAYER metal2 ;
  RECT 2554.180 0.000 2557.720 1.120 ;
  LAYER metal1 ;
  RECT 2554.180 0.000 2557.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2510.780 0.000 2514.320 1.120 ;
  LAYER metal4 ;
  RECT 2510.780 0.000 2514.320 1.120 ;
  LAYER metal3 ;
  RECT 2510.780 0.000 2514.320 1.120 ;
  LAYER metal2 ;
  RECT 2510.780 0.000 2514.320 1.120 ;
  LAYER metal1 ;
  RECT 2510.780 0.000 2514.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2502.100 0.000 2505.640 1.120 ;
  LAYER metal4 ;
  RECT 2502.100 0.000 2505.640 1.120 ;
  LAYER metal3 ;
  RECT 2502.100 0.000 2505.640 1.120 ;
  LAYER metal2 ;
  RECT 2502.100 0.000 2505.640 1.120 ;
  LAYER metal1 ;
  RECT 2502.100 0.000 2505.640 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2493.420 0.000 2496.960 1.120 ;
  LAYER metal4 ;
  RECT 2493.420 0.000 2496.960 1.120 ;
  LAYER metal3 ;
  RECT 2493.420 0.000 2496.960 1.120 ;
  LAYER metal2 ;
  RECT 2493.420 0.000 2496.960 1.120 ;
  LAYER metal1 ;
  RECT 2493.420 0.000 2496.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2484.740 0.000 2488.280 1.120 ;
  LAYER metal4 ;
  RECT 2484.740 0.000 2488.280 1.120 ;
  LAYER metal3 ;
  RECT 2484.740 0.000 2488.280 1.120 ;
  LAYER metal2 ;
  RECT 2484.740 0.000 2488.280 1.120 ;
  LAYER metal1 ;
  RECT 2484.740 0.000 2488.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2476.060 0.000 2479.600 1.120 ;
  LAYER metal4 ;
  RECT 2476.060 0.000 2479.600 1.120 ;
  LAYER metal3 ;
  RECT 2476.060 0.000 2479.600 1.120 ;
  LAYER metal2 ;
  RECT 2476.060 0.000 2479.600 1.120 ;
  LAYER metal1 ;
  RECT 2476.060 0.000 2479.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2467.380 0.000 2470.920 1.120 ;
  LAYER metal4 ;
  RECT 2467.380 0.000 2470.920 1.120 ;
  LAYER metal3 ;
  RECT 2467.380 0.000 2470.920 1.120 ;
  LAYER metal2 ;
  RECT 2467.380 0.000 2470.920 1.120 ;
  LAYER metal1 ;
  RECT 2467.380 0.000 2470.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2423.980 0.000 2427.520 1.120 ;
  LAYER metal4 ;
  RECT 2423.980 0.000 2427.520 1.120 ;
  LAYER metal3 ;
  RECT 2423.980 0.000 2427.520 1.120 ;
  LAYER metal2 ;
  RECT 2423.980 0.000 2427.520 1.120 ;
  LAYER metal1 ;
  RECT 2423.980 0.000 2427.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2415.300 0.000 2418.840 1.120 ;
  LAYER metal4 ;
  RECT 2415.300 0.000 2418.840 1.120 ;
  LAYER metal3 ;
  RECT 2415.300 0.000 2418.840 1.120 ;
  LAYER metal2 ;
  RECT 2415.300 0.000 2418.840 1.120 ;
  LAYER metal1 ;
  RECT 2415.300 0.000 2418.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2406.620 0.000 2410.160 1.120 ;
  LAYER metal4 ;
  RECT 2406.620 0.000 2410.160 1.120 ;
  LAYER metal3 ;
  RECT 2406.620 0.000 2410.160 1.120 ;
  LAYER metal2 ;
  RECT 2406.620 0.000 2410.160 1.120 ;
  LAYER metal1 ;
  RECT 2406.620 0.000 2410.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2397.940 0.000 2401.480 1.120 ;
  LAYER metal4 ;
  RECT 2397.940 0.000 2401.480 1.120 ;
  LAYER metal3 ;
  RECT 2397.940 0.000 2401.480 1.120 ;
  LAYER metal2 ;
  RECT 2397.940 0.000 2401.480 1.120 ;
  LAYER metal1 ;
  RECT 2397.940 0.000 2401.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2389.260 0.000 2392.800 1.120 ;
  LAYER metal4 ;
  RECT 2389.260 0.000 2392.800 1.120 ;
  LAYER metal3 ;
  RECT 2389.260 0.000 2392.800 1.120 ;
  LAYER metal2 ;
  RECT 2389.260 0.000 2392.800 1.120 ;
  LAYER metal1 ;
  RECT 2389.260 0.000 2392.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2380.580 0.000 2384.120 1.120 ;
  LAYER metal4 ;
  RECT 2380.580 0.000 2384.120 1.120 ;
  LAYER metal3 ;
  RECT 2380.580 0.000 2384.120 1.120 ;
  LAYER metal2 ;
  RECT 2380.580 0.000 2384.120 1.120 ;
  LAYER metal1 ;
  RECT 2380.580 0.000 2384.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2327.880 0.000 2331.420 1.120 ;
  LAYER metal4 ;
  RECT 2327.880 0.000 2331.420 1.120 ;
  LAYER metal3 ;
  RECT 2327.880 0.000 2331.420 1.120 ;
  LAYER metal2 ;
  RECT 2327.880 0.000 2331.420 1.120 ;
  LAYER metal1 ;
  RECT 2327.880 0.000 2331.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2314.240 0.000 2317.780 1.120 ;
  LAYER metal4 ;
  RECT 2314.240 0.000 2317.780 1.120 ;
  LAYER metal3 ;
  RECT 2314.240 0.000 2317.780 1.120 ;
  LAYER metal2 ;
  RECT 2314.240 0.000 2317.780 1.120 ;
  LAYER metal1 ;
  RECT 2314.240 0.000 2317.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2299.980 0.000 2303.520 1.120 ;
  LAYER metal4 ;
  RECT 2299.980 0.000 2303.520 1.120 ;
  LAYER metal3 ;
  RECT 2299.980 0.000 2303.520 1.120 ;
  LAYER metal2 ;
  RECT 2299.980 0.000 2303.520 1.120 ;
  LAYER metal1 ;
  RECT 2299.980 0.000 2303.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2291.300 0.000 2294.840 1.120 ;
  LAYER metal4 ;
  RECT 2291.300 0.000 2294.840 1.120 ;
  LAYER metal3 ;
  RECT 2291.300 0.000 2294.840 1.120 ;
  LAYER metal2 ;
  RECT 2291.300 0.000 2294.840 1.120 ;
  LAYER metal1 ;
  RECT 2291.300 0.000 2294.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2282.620 0.000 2286.160 1.120 ;
  LAYER metal4 ;
  RECT 2282.620 0.000 2286.160 1.120 ;
  LAYER metal3 ;
  RECT 2282.620 0.000 2286.160 1.120 ;
  LAYER metal2 ;
  RECT 2282.620 0.000 2286.160 1.120 ;
  LAYER metal1 ;
  RECT 2282.620 0.000 2286.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2273.940 0.000 2277.480 1.120 ;
  LAYER metal4 ;
  RECT 2273.940 0.000 2277.480 1.120 ;
  LAYER metal3 ;
  RECT 2273.940 0.000 2277.480 1.120 ;
  LAYER metal2 ;
  RECT 2273.940 0.000 2277.480 1.120 ;
  LAYER metal1 ;
  RECT 2273.940 0.000 2277.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2230.540 0.000 2234.080 1.120 ;
  LAYER metal4 ;
  RECT 2230.540 0.000 2234.080 1.120 ;
  LAYER metal3 ;
  RECT 2230.540 0.000 2234.080 1.120 ;
  LAYER metal2 ;
  RECT 2230.540 0.000 2234.080 1.120 ;
  LAYER metal1 ;
  RECT 2230.540 0.000 2234.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2221.860 0.000 2225.400 1.120 ;
  LAYER metal4 ;
  RECT 2221.860 0.000 2225.400 1.120 ;
  LAYER metal3 ;
  RECT 2221.860 0.000 2225.400 1.120 ;
  LAYER metal2 ;
  RECT 2221.860 0.000 2225.400 1.120 ;
  LAYER metal1 ;
  RECT 2221.860 0.000 2225.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2213.180 0.000 2216.720 1.120 ;
  LAYER metal4 ;
  RECT 2213.180 0.000 2216.720 1.120 ;
  LAYER metal3 ;
  RECT 2213.180 0.000 2216.720 1.120 ;
  LAYER metal2 ;
  RECT 2213.180 0.000 2216.720 1.120 ;
  LAYER metal1 ;
  RECT 2213.180 0.000 2216.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2204.500 0.000 2208.040 1.120 ;
  LAYER metal4 ;
  RECT 2204.500 0.000 2208.040 1.120 ;
  LAYER metal3 ;
  RECT 2204.500 0.000 2208.040 1.120 ;
  LAYER metal2 ;
  RECT 2204.500 0.000 2208.040 1.120 ;
  LAYER metal1 ;
  RECT 2204.500 0.000 2208.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2195.820 0.000 2199.360 1.120 ;
  LAYER metal4 ;
  RECT 2195.820 0.000 2199.360 1.120 ;
  LAYER metal3 ;
  RECT 2195.820 0.000 2199.360 1.120 ;
  LAYER metal2 ;
  RECT 2195.820 0.000 2199.360 1.120 ;
  LAYER metal1 ;
  RECT 2195.820 0.000 2199.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2187.140 0.000 2190.680 1.120 ;
  LAYER metal4 ;
  RECT 2187.140 0.000 2190.680 1.120 ;
  LAYER metal3 ;
  RECT 2187.140 0.000 2190.680 1.120 ;
  LAYER metal2 ;
  RECT 2187.140 0.000 2190.680 1.120 ;
  LAYER metal1 ;
  RECT 2187.140 0.000 2190.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2143.740 0.000 2147.280 1.120 ;
  LAYER metal4 ;
  RECT 2143.740 0.000 2147.280 1.120 ;
  LAYER metal3 ;
  RECT 2143.740 0.000 2147.280 1.120 ;
  LAYER metal2 ;
  RECT 2143.740 0.000 2147.280 1.120 ;
  LAYER metal1 ;
  RECT 2143.740 0.000 2147.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2135.060 0.000 2138.600 1.120 ;
  LAYER metal4 ;
  RECT 2135.060 0.000 2138.600 1.120 ;
  LAYER metal3 ;
  RECT 2135.060 0.000 2138.600 1.120 ;
  LAYER metal2 ;
  RECT 2135.060 0.000 2138.600 1.120 ;
  LAYER metal1 ;
  RECT 2135.060 0.000 2138.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2126.380 0.000 2129.920 1.120 ;
  LAYER metal4 ;
  RECT 2126.380 0.000 2129.920 1.120 ;
  LAYER metal3 ;
  RECT 2126.380 0.000 2129.920 1.120 ;
  LAYER metal2 ;
  RECT 2126.380 0.000 2129.920 1.120 ;
  LAYER metal1 ;
  RECT 2126.380 0.000 2129.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2117.700 0.000 2121.240 1.120 ;
  LAYER metal4 ;
  RECT 2117.700 0.000 2121.240 1.120 ;
  LAYER metal3 ;
  RECT 2117.700 0.000 2121.240 1.120 ;
  LAYER metal2 ;
  RECT 2117.700 0.000 2121.240 1.120 ;
  LAYER metal1 ;
  RECT 2117.700 0.000 2121.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2109.020 0.000 2112.560 1.120 ;
  LAYER metal4 ;
  RECT 2109.020 0.000 2112.560 1.120 ;
  LAYER metal3 ;
  RECT 2109.020 0.000 2112.560 1.120 ;
  LAYER metal2 ;
  RECT 2109.020 0.000 2112.560 1.120 ;
  LAYER metal1 ;
  RECT 2109.020 0.000 2112.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2100.340 0.000 2103.880 1.120 ;
  LAYER metal4 ;
  RECT 2100.340 0.000 2103.880 1.120 ;
  LAYER metal3 ;
  RECT 2100.340 0.000 2103.880 1.120 ;
  LAYER metal2 ;
  RECT 2100.340 0.000 2103.880 1.120 ;
  LAYER metal1 ;
  RECT 2100.340 0.000 2103.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2056.940 0.000 2060.480 1.120 ;
  LAYER metal4 ;
  RECT 2056.940 0.000 2060.480 1.120 ;
  LAYER metal3 ;
  RECT 2056.940 0.000 2060.480 1.120 ;
  LAYER metal2 ;
  RECT 2056.940 0.000 2060.480 1.120 ;
  LAYER metal1 ;
  RECT 2056.940 0.000 2060.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2048.260 0.000 2051.800 1.120 ;
  LAYER metal4 ;
  RECT 2048.260 0.000 2051.800 1.120 ;
  LAYER metal3 ;
  RECT 2048.260 0.000 2051.800 1.120 ;
  LAYER metal2 ;
  RECT 2048.260 0.000 2051.800 1.120 ;
  LAYER metal1 ;
  RECT 2048.260 0.000 2051.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2039.580 0.000 2043.120 1.120 ;
  LAYER metal4 ;
  RECT 2039.580 0.000 2043.120 1.120 ;
  LAYER metal3 ;
  RECT 2039.580 0.000 2043.120 1.120 ;
  LAYER metal2 ;
  RECT 2039.580 0.000 2043.120 1.120 ;
  LAYER metal1 ;
  RECT 2039.580 0.000 2043.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2030.900 0.000 2034.440 1.120 ;
  LAYER metal4 ;
  RECT 2030.900 0.000 2034.440 1.120 ;
  LAYER metal3 ;
  RECT 2030.900 0.000 2034.440 1.120 ;
  LAYER metal2 ;
  RECT 2030.900 0.000 2034.440 1.120 ;
  LAYER metal1 ;
  RECT 2030.900 0.000 2034.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2022.220 0.000 2025.760 1.120 ;
  LAYER metal4 ;
  RECT 2022.220 0.000 2025.760 1.120 ;
  LAYER metal3 ;
  RECT 2022.220 0.000 2025.760 1.120 ;
  LAYER metal2 ;
  RECT 2022.220 0.000 2025.760 1.120 ;
  LAYER metal1 ;
  RECT 2022.220 0.000 2025.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2013.540 0.000 2017.080 1.120 ;
  LAYER metal4 ;
  RECT 2013.540 0.000 2017.080 1.120 ;
  LAYER metal3 ;
  RECT 2013.540 0.000 2017.080 1.120 ;
  LAYER metal2 ;
  RECT 2013.540 0.000 2017.080 1.120 ;
  LAYER metal1 ;
  RECT 2013.540 0.000 2017.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1970.140 0.000 1973.680 1.120 ;
  LAYER metal4 ;
  RECT 1970.140 0.000 1973.680 1.120 ;
  LAYER metal3 ;
  RECT 1970.140 0.000 1973.680 1.120 ;
  LAYER metal2 ;
  RECT 1970.140 0.000 1973.680 1.120 ;
  LAYER metal1 ;
  RECT 1970.140 0.000 1973.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1961.460 0.000 1965.000 1.120 ;
  LAYER metal4 ;
  RECT 1961.460 0.000 1965.000 1.120 ;
  LAYER metal3 ;
  RECT 1961.460 0.000 1965.000 1.120 ;
  LAYER metal2 ;
  RECT 1961.460 0.000 1965.000 1.120 ;
  LAYER metal1 ;
  RECT 1961.460 0.000 1965.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1952.780 0.000 1956.320 1.120 ;
  LAYER metal4 ;
  RECT 1952.780 0.000 1956.320 1.120 ;
  LAYER metal3 ;
  RECT 1952.780 0.000 1956.320 1.120 ;
  LAYER metal2 ;
  RECT 1952.780 0.000 1956.320 1.120 ;
  LAYER metal1 ;
  RECT 1952.780 0.000 1956.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1944.100 0.000 1947.640 1.120 ;
  LAYER metal4 ;
  RECT 1944.100 0.000 1947.640 1.120 ;
  LAYER metal3 ;
  RECT 1944.100 0.000 1947.640 1.120 ;
  LAYER metal2 ;
  RECT 1944.100 0.000 1947.640 1.120 ;
  LAYER metal1 ;
  RECT 1944.100 0.000 1947.640 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1935.420 0.000 1938.960 1.120 ;
  LAYER metal4 ;
  RECT 1935.420 0.000 1938.960 1.120 ;
  LAYER metal3 ;
  RECT 1935.420 0.000 1938.960 1.120 ;
  LAYER metal2 ;
  RECT 1935.420 0.000 1938.960 1.120 ;
  LAYER metal1 ;
  RECT 1935.420 0.000 1938.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1926.740 0.000 1930.280 1.120 ;
  LAYER metal4 ;
  RECT 1926.740 0.000 1930.280 1.120 ;
  LAYER metal3 ;
  RECT 1926.740 0.000 1930.280 1.120 ;
  LAYER metal2 ;
  RECT 1926.740 0.000 1930.280 1.120 ;
  LAYER metal1 ;
  RECT 1926.740 0.000 1930.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1863.500 0.000 1867.040 1.120 ;
  LAYER metal4 ;
  RECT 1863.500 0.000 1867.040 1.120 ;
  LAYER metal3 ;
  RECT 1863.500 0.000 1867.040 1.120 ;
  LAYER metal2 ;
  RECT 1863.500 0.000 1867.040 1.120 ;
  LAYER metal1 ;
  RECT 1863.500 0.000 1867.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1854.820 0.000 1858.360 1.120 ;
  LAYER metal4 ;
  RECT 1854.820 0.000 1858.360 1.120 ;
  LAYER metal3 ;
  RECT 1854.820 0.000 1858.360 1.120 ;
  LAYER metal2 ;
  RECT 1854.820 0.000 1858.360 1.120 ;
  LAYER metal1 ;
  RECT 1854.820 0.000 1858.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1813.280 0.000 1816.820 1.120 ;
  LAYER metal4 ;
  RECT 1813.280 0.000 1816.820 1.120 ;
  LAYER metal3 ;
  RECT 1813.280 0.000 1816.820 1.120 ;
  LAYER metal2 ;
  RECT 1813.280 0.000 1816.820 1.120 ;
  LAYER metal1 ;
  RECT 1813.280 0.000 1816.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1789.100 0.000 1792.640 1.120 ;
  LAYER metal4 ;
  RECT 1789.100 0.000 1792.640 1.120 ;
  LAYER metal3 ;
  RECT 1789.100 0.000 1792.640 1.120 ;
  LAYER metal2 ;
  RECT 1789.100 0.000 1792.640 1.120 ;
  LAYER metal1 ;
  RECT 1789.100 0.000 1792.640 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1764.300 0.000 1767.840 1.120 ;
  LAYER metal4 ;
  RECT 1764.300 0.000 1767.840 1.120 ;
  LAYER metal3 ;
  RECT 1764.300 0.000 1767.840 1.120 ;
  LAYER metal2 ;
  RECT 1764.300 0.000 1767.840 1.120 ;
  LAYER metal1 ;
  RECT 1764.300 0.000 1767.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1738.260 0.000 1741.800 1.120 ;
  LAYER metal4 ;
  RECT 1738.260 0.000 1741.800 1.120 ;
  LAYER metal3 ;
  RECT 1738.260 0.000 1741.800 1.120 ;
  LAYER metal2 ;
  RECT 1738.260 0.000 1741.800 1.120 ;
  LAYER metal1 ;
  RECT 1738.260 0.000 1741.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1694.860 0.000 1698.400 1.120 ;
  LAYER metal4 ;
  RECT 1694.860 0.000 1698.400 1.120 ;
  LAYER metal3 ;
  RECT 1694.860 0.000 1698.400 1.120 ;
  LAYER metal2 ;
  RECT 1694.860 0.000 1698.400 1.120 ;
  LAYER metal1 ;
  RECT 1694.860 0.000 1698.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1686.180 0.000 1689.720 1.120 ;
  LAYER metal4 ;
  RECT 1686.180 0.000 1689.720 1.120 ;
  LAYER metal3 ;
  RECT 1686.180 0.000 1689.720 1.120 ;
  LAYER metal2 ;
  RECT 1686.180 0.000 1689.720 1.120 ;
  LAYER metal1 ;
  RECT 1686.180 0.000 1689.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1677.500 0.000 1681.040 1.120 ;
  LAYER metal4 ;
  RECT 1677.500 0.000 1681.040 1.120 ;
  LAYER metal3 ;
  RECT 1677.500 0.000 1681.040 1.120 ;
  LAYER metal2 ;
  RECT 1677.500 0.000 1681.040 1.120 ;
  LAYER metal1 ;
  RECT 1677.500 0.000 1681.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1668.820 0.000 1672.360 1.120 ;
  LAYER metal4 ;
  RECT 1668.820 0.000 1672.360 1.120 ;
  LAYER metal3 ;
  RECT 1668.820 0.000 1672.360 1.120 ;
  LAYER metal2 ;
  RECT 1668.820 0.000 1672.360 1.120 ;
  LAYER metal1 ;
  RECT 1668.820 0.000 1672.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1660.140 0.000 1663.680 1.120 ;
  LAYER metal4 ;
  RECT 1660.140 0.000 1663.680 1.120 ;
  LAYER metal3 ;
  RECT 1660.140 0.000 1663.680 1.120 ;
  LAYER metal2 ;
  RECT 1660.140 0.000 1663.680 1.120 ;
  LAYER metal1 ;
  RECT 1660.140 0.000 1663.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1651.460 0.000 1655.000 1.120 ;
  LAYER metal4 ;
  RECT 1651.460 0.000 1655.000 1.120 ;
  LAYER metal3 ;
  RECT 1651.460 0.000 1655.000 1.120 ;
  LAYER metal2 ;
  RECT 1651.460 0.000 1655.000 1.120 ;
  LAYER metal1 ;
  RECT 1651.460 0.000 1655.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1608.060 0.000 1611.600 1.120 ;
  LAYER metal4 ;
  RECT 1608.060 0.000 1611.600 1.120 ;
  LAYER metal3 ;
  RECT 1608.060 0.000 1611.600 1.120 ;
  LAYER metal2 ;
  RECT 1608.060 0.000 1611.600 1.120 ;
  LAYER metal1 ;
  RECT 1608.060 0.000 1611.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1599.380 0.000 1602.920 1.120 ;
  LAYER metal4 ;
  RECT 1599.380 0.000 1602.920 1.120 ;
  LAYER metal3 ;
  RECT 1599.380 0.000 1602.920 1.120 ;
  LAYER metal2 ;
  RECT 1599.380 0.000 1602.920 1.120 ;
  LAYER metal1 ;
  RECT 1599.380 0.000 1602.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1590.700 0.000 1594.240 1.120 ;
  LAYER metal4 ;
  RECT 1590.700 0.000 1594.240 1.120 ;
  LAYER metal3 ;
  RECT 1590.700 0.000 1594.240 1.120 ;
  LAYER metal2 ;
  RECT 1590.700 0.000 1594.240 1.120 ;
  LAYER metal1 ;
  RECT 1590.700 0.000 1594.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1582.020 0.000 1585.560 1.120 ;
  LAYER metal4 ;
  RECT 1582.020 0.000 1585.560 1.120 ;
  LAYER metal3 ;
  RECT 1582.020 0.000 1585.560 1.120 ;
  LAYER metal2 ;
  RECT 1582.020 0.000 1585.560 1.120 ;
  LAYER metal1 ;
  RECT 1582.020 0.000 1585.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1573.340 0.000 1576.880 1.120 ;
  LAYER metal4 ;
  RECT 1573.340 0.000 1576.880 1.120 ;
  LAYER metal3 ;
  RECT 1573.340 0.000 1576.880 1.120 ;
  LAYER metal2 ;
  RECT 1573.340 0.000 1576.880 1.120 ;
  LAYER metal1 ;
  RECT 1573.340 0.000 1576.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1564.660 0.000 1568.200 1.120 ;
  LAYER metal4 ;
  RECT 1564.660 0.000 1568.200 1.120 ;
  LAYER metal3 ;
  RECT 1564.660 0.000 1568.200 1.120 ;
  LAYER metal2 ;
  RECT 1564.660 0.000 1568.200 1.120 ;
  LAYER metal1 ;
  RECT 1564.660 0.000 1568.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1521.260 0.000 1524.800 1.120 ;
  LAYER metal4 ;
  RECT 1521.260 0.000 1524.800 1.120 ;
  LAYER metal3 ;
  RECT 1521.260 0.000 1524.800 1.120 ;
  LAYER metal2 ;
  RECT 1521.260 0.000 1524.800 1.120 ;
  LAYER metal1 ;
  RECT 1521.260 0.000 1524.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1512.580 0.000 1516.120 1.120 ;
  LAYER metal4 ;
  RECT 1512.580 0.000 1516.120 1.120 ;
  LAYER metal3 ;
  RECT 1512.580 0.000 1516.120 1.120 ;
  LAYER metal2 ;
  RECT 1512.580 0.000 1516.120 1.120 ;
  LAYER metal1 ;
  RECT 1512.580 0.000 1516.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1503.900 0.000 1507.440 1.120 ;
  LAYER metal4 ;
  RECT 1503.900 0.000 1507.440 1.120 ;
  LAYER metal3 ;
  RECT 1503.900 0.000 1507.440 1.120 ;
  LAYER metal2 ;
  RECT 1503.900 0.000 1507.440 1.120 ;
  LAYER metal1 ;
  RECT 1503.900 0.000 1507.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1495.220 0.000 1498.760 1.120 ;
  LAYER metal4 ;
  RECT 1495.220 0.000 1498.760 1.120 ;
  LAYER metal3 ;
  RECT 1495.220 0.000 1498.760 1.120 ;
  LAYER metal2 ;
  RECT 1495.220 0.000 1498.760 1.120 ;
  LAYER metal1 ;
  RECT 1495.220 0.000 1498.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1486.540 0.000 1490.080 1.120 ;
  LAYER metal4 ;
  RECT 1486.540 0.000 1490.080 1.120 ;
  LAYER metal3 ;
  RECT 1486.540 0.000 1490.080 1.120 ;
  LAYER metal2 ;
  RECT 1486.540 0.000 1490.080 1.120 ;
  LAYER metal1 ;
  RECT 1486.540 0.000 1490.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1477.860 0.000 1481.400 1.120 ;
  LAYER metal4 ;
  RECT 1477.860 0.000 1481.400 1.120 ;
  LAYER metal3 ;
  RECT 1477.860 0.000 1481.400 1.120 ;
  LAYER metal2 ;
  RECT 1477.860 0.000 1481.400 1.120 ;
  LAYER metal1 ;
  RECT 1477.860 0.000 1481.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1434.460 0.000 1438.000 1.120 ;
  LAYER metal4 ;
  RECT 1434.460 0.000 1438.000 1.120 ;
  LAYER metal3 ;
  RECT 1434.460 0.000 1438.000 1.120 ;
  LAYER metal2 ;
  RECT 1434.460 0.000 1438.000 1.120 ;
  LAYER metal1 ;
  RECT 1434.460 0.000 1438.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1425.780 0.000 1429.320 1.120 ;
  LAYER metal4 ;
  RECT 1425.780 0.000 1429.320 1.120 ;
  LAYER metal3 ;
  RECT 1425.780 0.000 1429.320 1.120 ;
  LAYER metal2 ;
  RECT 1425.780 0.000 1429.320 1.120 ;
  LAYER metal1 ;
  RECT 1425.780 0.000 1429.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1417.100 0.000 1420.640 1.120 ;
  LAYER metal4 ;
  RECT 1417.100 0.000 1420.640 1.120 ;
  LAYER metal3 ;
  RECT 1417.100 0.000 1420.640 1.120 ;
  LAYER metal2 ;
  RECT 1417.100 0.000 1420.640 1.120 ;
  LAYER metal1 ;
  RECT 1417.100 0.000 1420.640 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1408.420 0.000 1411.960 1.120 ;
  LAYER metal4 ;
  RECT 1408.420 0.000 1411.960 1.120 ;
  LAYER metal3 ;
  RECT 1408.420 0.000 1411.960 1.120 ;
  LAYER metal2 ;
  RECT 1408.420 0.000 1411.960 1.120 ;
  LAYER metal1 ;
  RECT 1408.420 0.000 1411.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1399.740 0.000 1403.280 1.120 ;
  LAYER metal4 ;
  RECT 1399.740 0.000 1403.280 1.120 ;
  LAYER metal3 ;
  RECT 1399.740 0.000 1403.280 1.120 ;
  LAYER metal2 ;
  RECT 1399.740 0.000 1403.280 1.120 ;
  LAYER metal1 ;
  RECT 1399.740 0.000 1403.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1391.060 0.000 1394.600 1.120 ;
  LAYER metal4 ;
  RECT 1391.060 0.000 1394.600 1.120 ;
  LAYER metal3 ;
  RECT 1391.060 0.000 1394.600 1.120 ;
  LAYER metal2 ;
  RECT 1391.060 0.000 1394.600 1.120 ;
  LAYER metal1 ;
  RECT 1391.060 0.000 1394.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1343.320 0.000 1346.860 1.120 ;
  LAYER metal4 ;
  RECT 1343.320 0.000 1346.860 1.120 ;
  LAYER metal3 ;
  RECT 1343.320 0.000 1346.860 1.120 ;
  LAYER metal2 ;
  RECT 1343.320 0.000 1346.860 1.120 ;
  LAYER metal1 ;
  RECT 1343.320 0.000 1346.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1329.680 0.000 1333.220 1.120 ;
  LAYER metal4 ;
  RECT 1329.680 0.000 1333.220 1.120 ;
  LAYER metal3 ;
  RECT 1329.680 0.000 1333.220 1.120 ;
  LAYER metal2 ;
  RECT 1329.680 0.000 1333.220 1.120 ;
  LAYER metal1 ;
  RECT 1329.680 0.000 1333.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1316.040 0.000 1319.580 1.120 ;
  LAYER metal4 ;
  RECT 1316.040 0.000 1319.580 1.120 ;
  LAYER metal3 ;
  RECT 1316.040 0.000 1319.580 1.120 ;
  LAYER metal2 ;
  RECT 1316.040 0.000 1319.580 1.120 ;
  LAYER metal1 ;
  RECT 1316.040 0.000 1319.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1301.780 0.000 1305.320 1.120 ;
  LAYER metal4 ;
  RECT 1301.780 0.000 1305.320 1.120 ;
  LAYER metal3 ;
  RECT 1301.780 0.000 1305.320 1.120 ;
  LAYER metal2 ;
  RECT 1301.780 0.000 1305.320 1.120 ;
  LAYER metal1 ;
  RECT 1301.780 0.000 1305.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1293.100 0.000 1296.640 1.120 ;
  LAYER metal4 ;
  RECT 1293.100 0.000 1296.640 1.120 ;
  LAYER metal3 ;
  RECT 1293.100 0.000 1296.640 1.120 ;
  LAYER metal2 ;
  RECT 1293.100 0.000 1296.640 1.120 ;
  LAYER metal1 ;
  RECT 1293.100 0.000 1296.640 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1284.420 0.000 1287.960 1.120 ;
  LAYER metal4 ;
  RECT 1284.420 0.000 1287.960 1.120 ;
  LAYER metal3 ;
  RECT 1284.420 0.000 1287.960 1.120 ;
  LAYER metal2 ;
  RECT 1284.420 0.000 1287.960 1.120 ;
  LAYER metal1 ;
  RECT 1284.420 0.000 1287.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1241.020 0.000 1244.560 1.120 ;
  LAYER metal4 ;
  RECT 1241.020 0.000 1244.560 1.120 ;
  LAYER metal3 ;
  RECT 1241.020 0.000 1244.560 1.120 ;
  LAYER metal2 ;
  RECT 1241.020 0.000 1244.560 1.120 ;
  LAYER metal1 ;
  RECT 1241.020 0.000 1244.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1232.340 0.000 1235.880 1.120 ;
  LAYER metal4 ;
  RECT 1232.340 0.000 1235.880 1.120 ;
  LAYER metal3 ;
  RECT 1232.340 0.000 1235.880 1.120 ;
  LAYER metal2 ;
  RECT 1232.340 0.000 1235.880 1.120 ;
  LAYER metal1 ;
  RECT 1232.340 0.000 1235.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1223.660 0.000 1227.200 1.120 ;
  LAYER metal4 ;
  RECT 1223.660 0.000 1227.200 1.120 ;
  LAYER metal3 ;
  RECT 1223.660 0.000 1227.200 1.120 ;
  LAYER metal2 ;
  RECT 1223.660 0.000 1227.200 1.120 ;
  LAYER metal1 ;
  RECT 1223.660 0.000 1227.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1214.980 0.000 1218.520 1.120 ;
  LAYER metal4 ;
  RECT 1214.980 0.000 1218.520 1.120 ;
  LAYER metal3 ;
  RECT 1214.980 0.000 1218.520 1.120 ;
  LAYER metal2 ;
  RECT 1214.980 0.000 1218.520 1.120 ;
  LAYER metal1 ;
  RECT 1214.980 0.000 1218.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1206.300 0.000 1209.840 1.120 ;
  LAYER metal4 ;
  RECT 1206.300 0.000 1209.840 1.120 ;
  LAYER metal3 ;
  RECT 1206.300 0.000 1209.840 1.120 ;
  LAYER metal2 ;
  RECT 1206.300 0.000 1209.840 1.120 ;
  LAYER metal1 ;
  RECT 1206.300 0.000 1209.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1197.620 0.000 1201.160 1.120 ;
  LAYER metal4 ;
  RECT 1197.620 0.000 1201.160 1.120 ;
  LAYER metal3 ;
  RECT 1197.620 0.000 1201.160 1.120 ;
  LAYER metal2 ;
  RECT 1197.620 0.000 1201.160 1.120 ;
  LAYER metal1 ;
  RECT 1197.620 0.000 1201.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1154.220 0.000 1157.760 1.120 ;
  LAYER metal4 ;
  RECT 1154.220 0.000 1157.760 1.120 ;
  LAYER metal3 ;
  RECT 1154.220 0.000 1157.760 1.120 ;
  LAYER metal2 ;
  RECT 1154.220 0.000 1157.760 1.120 ;
  LAYER metal1 ;
  RECT 1154.220 0.000 1157.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1145.540 0.000 1149.080 1.120 ;
  LAYER metal4 ;
  RECT 1145.540 0.000 1149.080 1.120 ;
  LAYER metal3 ;
  RECT 1145.540 0.000 1149.080 1.120 ;
  LAYER metal2 ;
  RECT 1145.540 0.000 1149.080 1.120 ;
  LAYER metal1 ;
  RECT 1145.540 0.000 1149.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1136.860 0.000 1140.400 1.120 ;
  LAYER metal4 ;
  RECT 1136.860 0.000 1140.400 1.120 ;
  LAYER metal3 ;
  RECT 1136.860 0.000 1140.400 1.120 ;
  LAYER metal2 ;
  RECT 1136.860 0.000 1140.400 1.120 ;
  LAYER metal1 ;
  RECT 1136.860 0.000 1140.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1128.180 0.000 1131.720 1.120 ;
  LAYER metal4 ;
  RECT 1128.180 0.000 1131.720 1.120 ;
  LAYER metal3 ;
  RECT 1128.180 0.000 1131.720 1.120 ;
  LAYER metal2 ;
  RECT 1128.180 0.000 1131.720 1.120 ;
  LAYER metal1 ;
  RECT 1128.180 0.000 1131.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1119.500 0.000 1123.040 1.120 ;
  LAYER metal4 ;
  RECT 1119.500 0.000 1123.040 1.120 ;
  LAYER metal3 ;
  RECT 1119.500 0.000 1123.040 1.120 ;
  LAYER metal2 ;
  RECT 1119.500 0.000 1123.040 1.120 ;
  LAYER metal1 ;
  RECT 1119.500 0.000 1123.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1110.820 0.000 1114.360 1.120 ;
  LAYER metal4 ;
  RECT 1110.820 0.000 1114.360 1.120 ;
  LAYER metal3 ;
  RECT 1110.820 0.000 1114.360 1.120 ;
  LAYER metal2 ;
  RECT 1110.820 0.000 1114.360 1.120 ;
  LAYER metal1 ;
  RECT 1110.820 0.000 1114.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1067.420 0.000 1070.960 1.120 ;
  LAYER metal4 ;
  RECT 1067.420 0.000 1070.960 1.120 ;
  LAYER metal3 ;
  RECT 1067.420 0.000 1070.960 1.120 ;
  LAYER metal2 ;
  RECT 1067.420 0.000 1070.960 1.120 ;
  LAYER metal1 ;
  RECT 1067.420 0.000 1070.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1058.740 0.000 1062.280 1.120 ;
  LAYER metal4 ;
  RECT 1058.740 0.000 1062.280 1.120 ;
  LAYER metal3 ;
  RECT 1058.740 0.000 1062.280 1.120 ;
  LAYER metal2 ;
  RECT 1058.740 0.000 1062.280 1.120 ;
  LAYER metal1 ;
  RECT 1058.740 0.000 1062.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1050.060 0.000 1053.600 1.120 ;
  LAYER metal4 ;
  RECT 1050.060 0.000 1053.600 1.120 ;
  LAYER metal3 ;
  RECT 1050.060 0.000 1053.600 1.120 ;
  LAYER metal2 ;
  RECT 1050.060 0.000 1053.600 1.120 ;
  LAYER metal1 ;
  RECT 1050.060 0.000 1053.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1041.380 0.000 1044.920 1.120 ;
  LAYER metal4 ;
  RECT 1041.380 0.000 1044.920 1.120 ;
  LAYER metal3 ;
  RECT 1041.380 0.000 1044.920 1.120 ;
  LAYER metal2 ;
  RECT 1041.380 0.000 1044.920 1.120 ;
  LAYER metal1 ;
  RECT 1041.380 0.000 1044.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1032.700 0.000 1036.240 1.120 ;
  LAYER metal4 ;
  RECT 1032.700 0.000 1036.240 1.120 ;
  LAYER metal3 ;
  RECT 1032.700 0.000 1036.240 1.120 ;
  LAYER metal2 ;
  RECT 1032.700 0.000 1036.240 1.120 ;
  LAYER metal1 ;
  RECT 1032.700 0.000 1036.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1024.020 0.000 1027.560 1.120 ;
  LAYER metal4 ;
  RECT 1024.020 0.000 1027.560 1.120 ;
  LAYER metal3 ;
  RECT 1024.020 0.000 1027.560 1.120 ;
  LAYER metal2 ;
  RECT 1024.020 0.000 1027.560 1.120 ;
  LAYER metal1 ;
  RECT 1024.020 0.000 1027.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 980.620 0.000 984.160 1.120 ;
  LAYER metal4 ;
  RECT 980.620 0.000 984.160 1.120 ;
  LAYER metal3 ;
  RECT 980.620 0.000 984.160 1.120 ;
  LAYER metal2 ;
  RECT 980.620 0.000 984.160 1.120 ;
  LAYER metal1 ;
  RECT 980.620 0.000 984.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 971.940 0.000 975.480 1.120 ;
  LAYER metal4 ;
  RECT 971.940 0.000 975.480 1.120 ;
  LAYER metal3 ;
  RECT 971.940 0.000 975.480 1.120 ;
  LAYER metal2 ;
  RECT 971.940 0.000 975.480 1.120 ;
  LAYER metal1 ;
  RECT 971.940 0.000 975.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 963.260 0.000 966.800 1.120 ;
  LAYER metal4 ;
  RECT 963.260 0.000 966.800 1.120 ;
  LAYER metal3 ;
  RECT 963.260 0.000 966.800 1.120 ;
  LAYER metal2 ;
  RECT 963.260 0.000 966.800 1.120 ;
  LAYER metal1 ;
  RECT 963.260 0.000 966.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 954.580 0.000 958.120 1.120 ;
  LAYER metal4 ;
  RECT 954.580 0.000 958.120 1.120 ;
  LAYER metal3 ;
  RECT 954.580 0.000 958.120 1.120 ;
  LAYER metal2 ;
  RECT 954.580 0.000 958.120 1.120 ;
  LAYER metal1 ;
  RECT 954.580 0.000 958.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 945.900 0.000 949.440 1.120 ;
  LAYER metal4 ;
  RECT 945.900 0.000 949.440 1.120 ;
  LAYER metal3 ;
  RECT 945.900 0.000 949.440 1.120 ;
  LAYER metal2 ;
  RECT 945.900 0.000 949.440 1.120 ;
  LAYER metal1 ;
  RECT 945.900 0.000 949.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 937.220 0.000 940.760 1.120 ;
  LAYER metal4 ;
  RECT 937.220 0.000 940.760 1.120 ;
  LAYER metal3 ;
  RECT 937.220 0.000 940.760 1.120 ;
  LAYER metal2 ;
  RECT 937.220 0.000 940.760 1.120 ;
  LAYER metal1 ;
  RECT 937.220 0.000 940.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 879.560 0.000 883.100 1.120 ;
  LAYER metal4 ;
  RECT 879.560 0.000 883.100 1.120 ;
  LAYER metal3 ;
  RECT 879.560 0.000 883.100 1.120 ;
  LAYER metal2 ;
  RECT 879.560 0.000 883.100 1.120 ;
  LAYER metal1 ;
  RECT 879.560 0.000 883.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 865.300 0.000 868.840 1.120 ;
  LAYER metal4 ;
  RECT 865.300 0.000 868.840 1.120 ;
  LAYER metal3 ;
  RECT 865.300 0.000 868.840 1.120 ;
  LAYER metal2 ;
  RECT 865.300 0.000 868.840 1.120 ;
  LAYER metal1 ;
  RECT 865.300 0.000 868.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 856.620 0.000 860.160 1.120 ;
  LAYER metal4 ;
  RECT 856.620 0.000 860.160 1.120 ;
  LAYER metal3 ;
  RECT 856.620 0.000 860.160 1.120 ;
  LAYER metal2 ;
  RECT 856.620 0.000 860.160 1.120 ;
  LAYER metal1 ;
  RECT 856.620 0.000 860.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 847.940 0.000 851.480 1.120 ;
  LAYER metal4 ;
  RECT 847.940 0.000 851.480 1.120 ;
  LAYER metal3 ;
  RECT 847.940 0.000 851.480 1.120 ;
  LAYER metal2 ;
  RECT 847.940 0.000 851.480 1.120 ;
  LAYER metal1 ;
  RECT 847.940 0.000 851.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 839.260 0.000 842.800 1.120 ;
  LAYER metal4 ;
  RECT 839.260 0.000 842.800 1.120 ;
  LAYER metal3 ;
  RECT 839.260 0.000 842.800 1.120 ;
  LAYER metal2 ;
  RECT 839.260 0.000 842.800 1.120 ;
  LAYER metal1 ;
  RECT 839.260 0.000 842.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 830.580 0.000 834.120 1.120 ;
  LAYER metal4 ;
  RECT 830.580 0.000 834.120 1.120 ;
  LAYER metal3 ;
  RECT 830.580 0.000 834.120 1.120 ;
  LAYER metal2 ;
  RECT 830.580 0.000 834.120 1.120 ;
  LAYER metal1 ;
  RECT 830.580 0.000 834.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 787.180 0.000 790.720 1.120 ;
  LAYER metal4 ;
  RECT 787.180 0.000 790.720 1.120 ;
  LAYER metal3 ;
  RECT 787.180 0.000 790.720 1.120 ;
  LAYER metal2 ;
  RECT 787.180 0.000 790.720 1.120 ;
  LAYER metal1 ;
  RECT 787.180 0.000 790.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 778.500 0.000 782.040 1.120 ;
  LAYER metal4 ;
  RECT 778.500 0.000 782.040 1.120 ;
  LAYER metal3 ;
  RECT 778.500 0.000 782.040 1.120 ;
  LAYER metal2 ;
  RECT 778.500 0.000 782.040 1.120 ;
  LAYER metal1 ;
  RECT 778.500 0.000 782.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 769.820 0.000 773.360 1.120 ;
  LAYER metal4 ;
  RECT 769.820 0.000 773.360 1.120 ;
  LAYER metal3 ;
  RECT 769.820 0.000 773.360 1.120 ;
  LAYER metal2 ;
  RECT 769.820 0.000 773.360 1.120 ;
  LAYER metal1 ;
  RECT 769.820 0.000 773.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 761.140 0.000 764.680 1.120 ;
  LAYER metal4 ;
  RECT 761.140 0.000 764.680 1.120 ;
  LAYER metal3 ;
  RECT 761.140 0.000 764.680 1.120 ;
  LAYER metal2 ;
  RECT 761.140 0.000 764.680 1.120 ;
  LAYER metal1 ;
  RECT 761.140 0.000 764.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 752.460 0.000 756.000 1.120 ;
  LAYER metal4 ;
  RECT 752.460 0.000 756.000 1.120 ;
  LAYER metal3 ;
  RECT 752.460 0.000 756.000 1.120 ;
  LAYER metal2 ;
  RECT 752.460 0.000 756.000 1.120 ;
  LAYER metal1 ;
  RECT 752.460 0.000 756.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 743.780 0.000 747.320 1.120 ;
  LAYER metal4 ;
  RECT 743.780 0.000 747.320 1.120 ;
  LAYER metal3 ;
  RECT 743.780 0.000 747.320 1.120 ;
  LAYER metal2 ;
  RECT 743.780 0.000 747.320 1.120 ;
  LAYER metal1 ;
  RECT 743.780 0.000 747.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 700.380 0.000 703.920 1.120 ;
  LAYER metal4 ;
  RECT 700.380 0.000 703.920 1.120 ;
  LAYER metal3 ;
  RECT 700.380 0.000 703.920 1.120 ;
  LAYER metal2 ;
  RECT 700.380 0.000 703.920 1.120 ;
  LAYER metal1 ;
  RECT 700.380 0.000 703.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 691.700 0.000 695.240 1.120 ;
  LAYER metal4 ;
  RECT 691.700 0.000 695.240 1.120 ;
  LAYER metal3 ;
  RECT 691.700 0.000 695.240 1.120 ;
  LAYER metal2 ;
  RECT 691.700 0.000 695.240 1.120 ;
  LAYER metal1 ;
  RECT 691.700 0.000 695.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 683.020 0.000 686.560 1.120 ;
  LAYER metal4 ;
  RECT 683.020 0.000 686.560 1.120 ;
  LAYER metal3 ;
  RECT 683.020 0.000 686.560 1.120 ;
  LAYER metal2 ;
  RECT 683.020 0.000 686.560 1.120 ;
  LAYER metal1 ;
  RECT 683.020 0.000 686.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 674.340 0.000 677.880 1.120 ;
  LAYER metal4 ;
  RECT 674.340 0.000 677.880 1.120 ;
  LAYER metal3 ;
  RECT 674.340 0.000 677.880 1.120 ;
  LAYER metal2 ;
  RECT 674.340 0.000 677.880 1.120 ;
  LAYER metal1 ;
  RECT 674.340 0.000 677.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 665.660 0.000 669.200 1.120 ;
  LAYER metal4 ;
  RECT 665.660 0.000 669.200 1.120 ;
  LAYER metal3 ;
  RECT 665.660 0.000 669.200 1.120 ;
  LAYER metal2 ;
  RECT 665.660 0.000 669.200 1.120 ;
  LAYER metal1 ;
  RECT 665.660 0.000 669.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 656.980 0.000 660.520 1.120 ;
  LAYER metal4 ;
  RECT 656.980 0.000 660.520 1.120 ;
  LAYER metal3 ;
  RECT 656.980 0.000 660.520 1.120 ;
  LAYER metal2 ;
  RECT 656.980 0.000 660.520 1.120 ;
  LAYER metal1 ;
  RECT 656.980 0.000 660.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 613.580 0.000 617.120 1.120 ;
  LAYER metal4 ;
  RECT 613.580 0.000 617.120 1.120 ;
  LAYER metal3 ;
  RECT 613.580 0.000 617.120 1.120 ;
  LAYER metal2 ;
  RECT 613.580 0.000 617.120 1.120 ;
  LAYER metal1 ;
  RECT 613.580 0.000 617.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 604.900 0.000 608.440 1.120 ;
  LAYER metal4 ;
  RECT 604.900 0.000 608.440 1.120 ;
  LAYER metal3 ;
  RECT 604.900 0.000 608.440 1.120 ;
  LAYER metal2 ;
  RECT 604.900 0.000 608.440 1.120 ;
  LAYER metal1 ;
  RECT 604.900 0.000 608.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 596.220 0.000 599.760 1.120 ;
  LAYER metal4 ;
  RECT 596.220 0.000 599.760 1.120 ;
  LAYER metal3 ;
  RECT 596.220 0.000 599.760 1.120 ;
  LAYER metal2 ;
  RECT 596.220 0.000 599.760 1.120 ;
  LAYER metal1 ;
  RECT 596.220 0.000 599.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 587.540 0.000 591.080 1.120 ;
  LAYER metal4 ;
  RECT 587.540 0.000 591.080 1.120 ;
  LAYER metal3 ;
  RECT 587.540 0.000 591.080 1.120 ;
  LAYER metal2 ;
  RECT 587.540 0.000 591.080 1.120 ;
  LAYER metal1 ;
  RECT 587.540 0.000 591.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 578.860 0.000 582.400 1.120 ;
  LAYER metal4 ;
  RECT 578.860 0.000 582.400 1.120 ;
  LAYER metal3 ;
  RECT 578.860 0.000 582.400 1.120 ;
  LAYER metal2 ;
  RECT 578.860 0.000 582.400 1.120 ;
  LAYER metal1 ;
  RECT 578.860 0.000 582.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal4 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal3 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal2 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal1 ;
  RECT 570.180 0.000 573.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 526.780 0.000 530.320 1.120 ;
  LAYER metal4 ;
  RECT 526.780 0.000 530.320 1.120 ;
  LAYER metal3 ;
  RECT 526.780 0.000 530.320 1.120 ;
  LAYER metal2 ;
  RECT 526.780 0.000 530.320 1.120 ;
  LAYER metal1 ;
  RECT 526.780 0.000 530.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 518.100 0.000 521.640 1.120 ;
  LAYER metal4 ;
  RECT 518.100 0.000 521.640 1.120 ;
  LAYER metal3 ;
  RECT 518.100 0.000 521.640 1.120 ;
  LAYER metal2 ;
  RECT 518.100 0.000 521.640 1.120 ;
  LAYER metal1 ;
  RECT 518.100 0.000 521.640 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 509.420 0.000 512.960 1.120 ;
  LAYER metal4 ;
  RECT 509.420 0.000 512.960 1.120 ;
  LAYER metal3 ;
  RECT 509.420 0.000 512.960 1.120 ;
  LAYER metal2 ;
  RECT 509.420 0.000 512.960 1.120 ;
  LAYER metal1 ;
  RECT 509.420 0.000 512.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 500.740 0.000 504.280 1.120 ;
  LAYER metal4 ;
  RECT 500.740 0.000 504.280 1.120 ;
  LAYER metal3 ;
  RECT 500.740 0.000 504.280 1.120 ;
  LAYER metal2 ;
  RECT 500.740 0.000 504.280 1.120 ;
  LAYER metal1 ;
  RECT 500.740 0.000 504.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 492.060 0.000 495.600 1.120 ;
  LAYER metal4 ;
  RECT 492.060 0.000 495.600 1.120 ;
  LAYER metal3 ;
  RECT 492.060 0.000 495.600 1.120 ;
  LAYER metal2 ;
  RECT 492.060 0.000 495.600 1.120 ;
  LAYER metal1 ;
  RECT 492.060 0.000 495.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 478.420 0.000 481.960 1.120 ;
  LAYER metal4 ;
  RECT 478.420 0.000 481.960 1.120 ;
  LAYER metal3 ;
  RECT 478.420 0.000 481.960 1.120 ;
  LAYER metal2 ;
  RECT 478.420 0.000 481.960 1.120 ;
  LAYER metal1 ;
  RECT 478.420 0.000 481.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 419.520 0.000 423.060 1.120 ;
  LAYER metal4 ;
  RECT 419.520 0.000 423.060 1.120 ;
  LAYER metal3 ;
  RECT 419.520 0.000 423.060 1.120 ;
  LAYER metal2 ;
  RECT 419.520 0.000 423.060 1.120 ;
  LAYER metal1 ;
  RECT 419.520 0.000 423.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 410.840 0.000 414.380 1.120 ;
  LAYER metal4 ;
  RECT 410.840 0.000 414.380 1.120 ;
  LAYER metal3 ;
  RECT 410.840 0.000 414.380 1.120 ;
  LAYER metal2 ;
  RECT 410.840 0.000 414.380 1.120 ;
  LAYER metal1 ;
  RECT 410.840 0.000 414.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 402.160 0.000 405.700 1.120 ;
  LAYER metal4 ;
  RECT 402.160 0.000 405.700 1.120 ;
  LAYER metal3 ;
  RECT 402.160 0.000 405.700 1.120 ;
  LAYER metal2 ;
  RECT 402.160 0.000 405.700 1.120 ;
  LAYER metal1 ;
  RECT 402.160 0.000 405.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 393.480 0.000 397.020 1.120 ;
  LAYER metal4 ;
  RECT 393.480 0.000 397.020 1.120 ;
  LAYER metal3 ;
  RECT 393.480 0.000 397.020 1.120 ;
  LAYER metal2 ;
  RECT 393.480 0.000 397.020 1.120 ;
  LAYER metal1 ;
  RECT 393.480 0.000 397.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 384.800 0.000 388.340 1.120 ;
  LAYER metal4 ;
  RECT 384.800 0.000 388.340 1.120 ;
  LAYER metal3 ;
  RECT 384.800 0.000 388.340 1.120 ;
  LAYER metal2 ;
  RECT 384.800 0.000 388.340 1.120 ;
  LAYER metal1 ;
  RECT 384.800 0.000 388.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 376.120 0.000 379.660 1.120 ;
  LAYER metal4 ;
  RECT 376.120 0.000 379.660 1.120 ;
  LAYER metal3 ;
  RECT 376.120 0.000 379.660 1.120 ;
  LAYER metal2 ;
  RECT 376.120 0.000 379.660 1.120 ;
  LAYER metal1 ;
  RECT 376.120 0.000 379.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 332.720 0.000 336.260 1.120 ;
  LAYER metal4 ;
  RECT 332.720 0.000 336.260 1.120 ;
  LAYER metal3 ;
  RECT 332.720 0.000 336.260 1.120 ;
  LAYER metal2 ;
  RECT 332.720 0.000 336.260 1.120 ;
  LAYER metal1 ;
  RECT 332.720 0.000 336.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 324.040 0.000 327.580 1.120 ;
  LAYER metal4 ;
  RECT 324.040 0.000 327.580 1.120 ;
  LAYER metal3 ;
  RECT 324.040 0.000 327.580 1.120 ;
  LAYER metal2 ;
  RECT 324.040 0.000 327.580 1.120 ;
  LAYER metal1 ;
  RECT 324.040 0.000 327.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 315.360 0.000 318.900 1.120 ;
  LAYER metal4 ;
  RECT 315.360 0.000 318.900 1.120 ;
  LAYER metal3 ;
  RECT 315.360 0.000 318.900 1.120 ;
  LAYER metal2 ;
  RECT 315.360 0.000 318.900 1.120 ;
  LAYER metal1 ;
  RECT 315.360 0.000 318.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 306.680 0.000 310.220 1.120 ;
  LAYER metal4 ;
  RECT 306.680 0.000 310.220 1.120 ;
  LAYER metal3 ;
  RECT 306.680 0.000 310.220 1.120 ;
  LAYER metal2 ;
  RECT 306.680 0.000 310.220 1.120 ;
  LAYER metal1 ;
  RECT 306.680 0.000 310.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 298.000 0.000 301.540 1.120 ;
  LAYER metal4 ;
  RECT 298.000 0.000 301.540 1.120 ;
  LAYER metal3 ;
  RECT 298.000 0.000 301.540 1.120 ;
  LAYER metal2 ;
  RECT 298.000 0.000 301.540 1.120 ;
  LAYER metal1 ;
  RECT 298.000 0.000 301.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 289.320 0.000 292.860 1.120 ;
  LAYER metal4 ;
  RECT 289.320 0.000 292.860 1.120 ;
  LAYER metal3 ;
  RECT 289.320 0.000 292.860 1.120 ;
  LAYER metal2 ;
  RECT 289.320 0.000 292.860 1.120 ;
  LAYER metal1 ;
  RECT 289.320 0.000 292.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 245.920 0.000 249.460 1.120 ;
  LAYER metal4 ;
  RECT 245.920 0.000 249.460 1.120 ;
  LAYER metal3 ;
  RECT 245.920 0.000 249.460 1.120 ;
  LAYER metal2 ;
  RECT 245.920 0.000 249.460 1.120 ;
  LAYER metal1 ;
  RECT 245.920 0.000 249.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 237.240 0.000 240.780 1.120 ;
  LAYER metal4 ;
  RECT 237.240 0.000 240.780 1.120 ;
  LAYER metal3 ;
  RECT 237.240 0.000 240.780 1.120 ;
  LAYER metal2 ;
  RECT 237.240 0.000 240.780 1.120 ;
  LAYER metal1 ;
  RECT 237.240 0.000 240.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 228.560 0.000 232.100 1.120 ;
  LAYER metal4 ;
  RECT 228.560 0.000 232.100 1.120 ;
  LAYER metal3 ;
  RECT 228.560 0.000 232.100 1.120 ;
  LAYER metal2 ;
  RECT 228.560 0.000 232.100 1.120 ;
  LAYER metal1 ;
  RECT 228.560 0.000 232.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 219.880 0.000 223.420 1.120 ;
  LAYER metal4 ;
  RECT 219.880 0.000 223.420 1.120 ;
  LAYER metal3 ;
  RECT 219.880 0.000 223.420 1.120 ;
  LAYER metal2 ;
  RECT 219.880 0.000 223.420 1.120 ;
  LAYER metal1 ;
  RECT 219.880 0.000 223.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 211.200 0.000 214.740 1.120 ;
  LAYER metal4 ;
  RECT 211.200 0.000 214.740 1.120 ;
  LAYER metal3 ;
  RECT 211.200 0.000 214.740 1.120 ;
  LAYER metal2 ;
  RECT 211.200 0.000 214.740 1.120 ;
  LAYER metal1 ;
  RECT 211.200 0.000 214.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 202.520 0.000 206.060 1.120 ;
  LAYER metal4 ;
  RECT 202.520 0.000 206.060 1.120 ;
  LAYER metal3 ;
  RECT 202.520 0.000 206.060 1.120 ;
  LAYER metal2 ;
  RECT 202.520 0.000 206.060 1.120 ;
  LAYER metal1 ;
  RECT 202.520 0.000 206.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 159.120 0.000 162.660 1.120 ;
  LAYER metal4 ;
  RECT 159.120 0.000 162.660 1.120 ;
  LAYER metal3 ;
  RECT 159.120 0.000 162.660 1.120 ;
  LAYER metal2 ;
  RECT 159.120 0.000 162.660 1.120 ;
  LAYER metal1 ;
  RECT 159.120 0.000 162.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 150.440 0.000 153.980 1.120 ;
  LAYER metal4 ;
  RECT 150.440 0.000 153.980 1.120 ;
  LAYER metal3 ;
  RECT 150.440 0.000 153.980 1.120 ;
  LAYER metal2 ;
  RECT 150.440 0.000 153.980 1.120 ;
  LAYER metal1 ;
  RECT 150.440 0.000 153.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 141.760 0.000 145.300 1.120 ;
  LAYER metal4 ;
  RECT 141.760 0.000 145.300 1.120 ;
  LAYER metal3 ;
  RECT 141.760 0.000 145.300 1.120 ;
  LAYER metal2 ;
  RECT 141.760 0.000 145.300 1.120 ;
  LAYER metal1 ;
  RECT 141.760 0.000 145.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 133.080 0.000 136.620 1.120 ;
  LAYER metal4 ;
  RECT 133.080 0.000 136.620 1.120 ;
  LAYER metal3 ;
  RECT 133.080 0.000 136.620 1.120 ;
  LAYER metal2 ;
  RECT 133.080 0.000 136.620 1.120 ;
  LAYER metal1 ;
  RECT 133.080 0.000 136.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 124.400 0.000 127.940 1.120 ;
  LAYER metal4 ;
  RECT 124.400 0.000 127.940 1.120 ;
  LAYER metal3 ;
  RECT 124.400 0.000 127.940 1.120 ;
  LAYER metal2 ;
  RECT 124.400 0.000 127.940 1.120 ;
  LAYER metal1 ;
  RECT 124.400 0.000 127.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 115.720 0.000 119.260 1.120 ;
  LAYER metal4 ;
  RECT 115.720 0.000 119.260 1.120 ;
  LAYER metal3 ;
  RECT 115.720 0.000 119.260 1.120 ;
  LAYER metal2 ;
  RECT 115.720 0.000 119.260 1.120 ;
  LAYER metal1 ;
  RECT 115.720 0.000 119.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 72.320 0.000 75.860 1.120 ;
  LAYER metal4 ;
  RECT 72.320 0.000 75.860 1.120 ;
  LAYER metal3 ;
  RECT 72.320 0.000 75.860 1.120 ;
  LAYER metal2 ;
  RECT 72.320 0.000 75.860 1.120 ;
  LAYER metal1 ;
  RECT 72.320 0.000 75.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 63.640 0.000 67.180 1.120 ;
  LAYER metal4 ;
  RECT 63.640 0.000 67.180 1.120 ;
  LAYER metal3 ;
  RECT 63.640 0.000 67.180 1.120 ;
  LAYER metal2 ;
  RECT 63.640 0.000 67.180 1.120 ;
  LAYER metal1 ;
  RECT 63.640 0.000 67.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER metal4 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER metal3 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER metal2 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER metal1 ;
  RECT 54.960 0.000 58.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER metal4 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER metal3 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER metal2 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER metal1 ;
  RECT 41.940 0.000 45.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER metal4 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER metal3 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER metal2 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER metal1 ;
  RECT 28.300 0.000 31.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 14.660 0.000 18.200 1.120 ;
  LAYER metal4 ;
  RECT 14.660 0.000 18.200 1.120 ;
  LAYER metal3 ;
  RECT 14.660 0.000 18.200 1.120 ;
  LAYER metal2 ;
  RECT 14.660 0.000 18.200 1.120 ;
  LAYER metal1 ;
  RECT 14.660 0.000 18.200 1.120 ;
 END
END GND
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal5 ;
  RECT 3612.860 1693.220 3613.980 1696.460 ;
  LAYER metal4 ;
  RECT 3612.860 1693.220 3613.980 1696.460 ;
  LAYER metal3 ;
  RECT 3612.860 1693.220 3613.980 1696.460 ;
  LAYER metal2 ;
  RECT 3612.860 1693.220 3613.980 1696.460 ;
  LAYER metal1 ;
  RECT 3612.860 1693.220 3613.980 1696.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1685.380 3613.980 1688.620 ;
  LAYER metal4 ;
  RECT 3612.860 1685.380 3613.980 1688.620 ;
  LAYER metal3 ;
  RECT 3612.860 1685.380 3613.980 1688.620 ;
  LAYER metal2 ;
  RECT 3612.860 1685.380 3613.980 1688.620 ;
  LAYER metal1 ;
  RECT 3612.860 1685.380 3613.980 1688.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1677.540 3613.980 1680.780 ;
  LAYER metal4 ;
  RECT 3612.860 1677.540 3613.980 1680.780 ;
  LAYER metal3 ;
  RECT 3612.860 1677.540 3613.980 1680.780 ;
  LAYER metal2 ;
  RECT 3612.860 1677.540 3613.980 1680.780 ;
  LAYER metal1 ;
  RECT 3612.860 1677.540 3613.980 1680.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1669.700 3613.980 1672.940 ;
  LAYER metal4 ;
  RECT 3612.860 1669.700 3613.980 1672.940 ;
  LAYER metal3 ;
  RECT 3612.860 1669.700 3613.980 1672.940 ;
  LAYER metal2 ;
  RECT 3612.860 1669.700 3613.980 1672.940 ;
  LAYER metal1 ;
  RECT 3612.860 1669.700 3613.980 1672.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1661.860 3613.980 1665.100 ;
  LAYER metal4 ;
  RECT 3612.860 1661.860 3613.980 1665.100 ;
  LAYER metal3 ;
  RECT 3612.860 1661.860 3613.980 1665.100 ;
  LAYER metal2 ;
  RECT 3612.860 1661.860 3613.980 1665.100 ;
  LAYER metal1 ;
  RECT 3612.860 1661.860 3613.980 1665.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1654.020 3613.980 1657.260 ;
  LAYER metal4 ;
  RECT 3612.860 1654.020 3613.980 1657.260 ;
  LAYER metal3 ;
  RECT 3612.860 1654.020 3613.980 1657.260 ;
  LAYER metal2 ;
  RECT 3612.860 1654.020 3613.980 1657.260 ;
  LAYER metal1 ;
  RECT 3612.860 1654.020 3613.980 1657.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1614.820 3613.980 1618.060 ;
  LAYER metal4 ;
  RECT 3612.860 1614.820 3613.980 1618.060 ;
  LAYER metal3 ;
  RECT 3612.860 1614.820 3613.980 1618.060 ;
  LAYER metal2 ;
  RECT 3612.860 1614.820 3613.980 1618.060 ;
  LAYER metal1 ;
  RECT 3612.860 1614.820 3613.980 1618.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1606.980 3613.980 1610.220 ;
  LAYER metal4 ;
  RECT 3612.860 1606.980 3613.980 1610.220 ;
  LAYER metal3 ;
  RECT 3612.860 1606.980 3613.980 1610.220 ;
  LAYER metal2 ;
  RECT 3612.860 1606.980 3613.980 1610.220 ;
  LAYER metal1 ;
  RECT 3612.860 1606.980 3613.980 1610.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1599.140 3613.980 1602.380 ;
  LAYER metal4 ;
  RECT 3612.860 1599.140 3613.980 1602.380 ;
  LAYER metal3 ;
  RECT 3612.860 1599.140 3613.980 1602.380 ;
  LAYER metal2 ;
  RECT 3612.860 1599.140 3613.980 1602.380 ;
  LAYER metal1 ;
  RECT 3612.860 1599.140 3613.980 1602.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1591.300 3613.980 1594.540 ;
  LAYER metal4 ;
  RECT 3612.860 1591.300 3613.980 1594.540 ;
  LAYER metal3 ;
  RECT 3612.860 1591.300 3613.980 1594.540 ;
  LAYER metal2 ;
  RECT 3612.860 1591.300 3613.980 1594.540 ;
  LAYER metal1 ;
  RECT 3612.860 1591.300 3613.980 1594.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1583.460 3613.980 1586.700 ;
  LAYER metal4 ;
  RECT 3612.860 1583.460 3613.980 1586.700 ;
  LAYER metal3 ;
  RECT 3612.860 1583.460 3613.980 1586.700 ;
  LAYER metal2 ;
  RECT 3612.860 1583.460 3613.980 1586.700 ;
  LAYER metal1 ;
  RECT 3612.860 1583.460 3613.980 1586.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1575.620 3613.980 1578.860 ;
  LAYER metal4 ;
  RECT 3612.860 1575.620 3613.980 1578.860 ;
  LAYER metal3 ;
  RECT 3612.860 1575.620 3613.980 1578.860 ;
  LAYER metal2 ;
  RECT 3612.860 1575.620 3613.980 1578.860 ;
  LAYER metal1 ;
  RECT 3612.860 1575.620 3613.980 1578.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1536.420 3613.980 1539.660 ;
  LAYER metal4 ;
  RECT 3612.860 1536.420 3613.980 1539.660 ;
  LAYER metal3 ;
  RECT 3612.860 1536.420 3613.980 1539.660 ;
  LAYER metal2 ;
  RECT 3612.860 1536.420 3613.980 1539.660 ;
  LAYER metal1 ;
  RECT 3612.860 1536.420 3613.980 1539.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1528.580 3613.980 1531.820 ;
  LAYER metal4 ;
  RECT 3612.860 1528.580 3613.980 1531.820 ;
  LAYER metal3 ;
  RECT 3612.860 1528.580 3613.980 1531.820 ;
  LAYER metal2 ;
  RECT 3612.860 1528.580 3613.980 1531.820 ;
  LAYER metal1 ;
  RECT 3612.860 1528.580 3613.980 1531.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1520.740 3613.980 1523.980 ;
  LAYER metal4 ;
  RECT 3612.860 1520.740 3613.980 1523.980 ;
  LAYER metal3 ;
  RECT 3612.860 1520.740 3613.980 1523.980 ;
  LAYER metal2 ;
  RECT 3612.860 1520.740 3613.980 1523.980 ;
  LAYER metal1 ;
  RECT 3612.860 1520.740 3613.980 1523.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1512.900 3613.980 1516.140 ;
  LAYER metal4 ;
  RECT 3612.860 1512.900 3613.980 1516.140 ;
  LAYER metal3 ;
  RECT 3612.860 1512.900 3613.980 1516.140 ;
  LAYER metal2 ;
  RECT 3612.860 1512.900 3613.980 1516.140 ;
  LAYER metal1 ;
  RECT 3612.860 1512.900 3613.980 1516.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1505.060 3613.980 1508.300 ;
  LAYER metal4 ;
  RECT 3612.860 1505.060 3613.980 1508.300 ;
  LAYER metal3 ;
  RECT 3612.860 1505.060 3613.980 1508.300 ;
  LAYER metal2 ;
  RECT 3612.860 1505.060 3613.980 1508.300 ;
  LAYER metal1 ;
  RECT 3612.860 1505.060 3613.980 1508.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1497.220 3613.980 1500.460 ;
  LAYER metal4 ;
  RECT 3612.860 1497.220 3613.980 1500.460 ;
  LAYER metal3 ;
  RECT 3612.860 1497.220 3613.980 1500.460 ;
  LAYER metal2 ;
  RECT 3612.860 1497.220 3613.980 1500.460 ;
  LAYER metal1 ;
  RECT 3612.860 1497.220 3613.980 1500.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1458.020 3613.980 1461.260 ;
  LAYER metal4 ;
  RECT 3612.860 1458.020 3613.980 1461.260 ;
  LAYER metal3 ;
  RECT 3612.860 1458.020 3613.980 1461.260 ;
  LAYER metal2 ;
  RECT 3612.860 1458.020 3613.980 1461.260 ;
  LAYER metal1 ;
  RECT 3612.860 1458.020 3613.980 1461.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1450.180 3613.980 1453.420 ;
  LAYER metal4 ;
  RECT 3612.860 1450.180 3613.980 1453.420 ;
  LAYER metal3 ;
  RECT 3612.860 1450.180 3613.980 1453.420 ;
  LAYER metal2 ;
  RECT 3612.860 1450.180 3613.980 1453.420 ;
  LAYER metal1 ;
  RECT 3612.860 1450.180 3613.980 1453.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1442.340 3613.980 1445.580 ;
  LAYER metal4 ;
  RECT 3612.860 1442.340 3613.980 1445.580 ;
  LAYER metal3 ;
  RECT 3612.860 1442.340 3613.980 1445.580 ;
  LAYER metal2 ;
  RECT 3612.860 1442.340 3613.980 1445.580 ;
  LAYER metal1 ;
  RECT 3612.860 1442.340 3613.980 1445.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1434.500 3613.980 1437.740 ;
  LAYER metal4 ;
  RECT 3612.860 1434.500 3613.980 1437.740 ;
  LAYER metal3 ;
  RECT 3612.860 1434.500 3613.980 1437.740 ;
  LAYER metal2 ;
  RECT 3612.860 1434.500 3613.980 1437.740 ;
  LAYER metal1 ;
  RECT 3612.860 1434.500 3613.980 1437.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1426.660 3613.980 1429.900 ;
  LAYER metal4 ;
  RECT 3612.860 1426.660 3613.980 1429.900 ;
  LAYER metal3 ;
  RECT 3612.860 1426.660 3613.980 1429.900 ;
  LAYER metal2 ;
  RECT 3612.860 1426.660 3613.980 1429.900 ;
  LAYER metal1 ;
  RECT 3612.860 1426.660 3613.980 1429.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1418.820 3613.980 1422.060 ;
  LAYER metal4 ;
  RECT 3612.860 1418.820 3613.980 1422.060 ;
  LAYER metal3 ;
  RECT 3612.860 1418.820 3613.980 1422.060 ;
  LAYER metal2 ;
  RECT 3612.860 1418.820 3613.980 1422.060 ;
  LAYER metal1 ;
  RECT 3612.860 1418.820 3613.980 1422.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1379.620 3613.980 1382.860 ;
  LAYER metal4 ;
  RECT 3612.860 1379.620 3613.980 1382.860 ;
  LAYER metal3 ;
  RECT 3612.860 1379.620 3613.980 1382.860 ;
  LAYER metal2 ;
  RECT 3612.860 1379.620 3613.980 1382.860 ;
  LAYER metal1 ;
  RECT 3612.860 1379.620 3613.980 1382.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1371.780 3613.980 1375.020 ;
  LAYER metal4 ;
  RECT 3612.860 1371.780 3613.980 1375.020 ;
  LAYER metal3 ;
  RECT 3612.860 1371.780 3613.980 1375.020 ;
  LAYER metal2 ;
  RECT 3612.860 1371.780 3613.980 1375.020 ;
  LAYER metal1 ;
  RECT 3612.860 1371.780 3613.980 1375.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1363.940 3613.980 1367.180 ;
  LAYER metal4 ;
  RECT 3612.860 1363.940 3613.980 1367.180 ;
  LAYER metal3 ;
  RECT 3612.860 1363.940 3613.980 1367.180 ;
  LAYER metal2 ;
  RECT 3612.860 1363.940 3613.980 1367.180 ;
  LAYER metal1 ;
  RECT 3612.860 1363.940 3613.980 1367.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1356.100 3613.980 1359.340 ;
  LAYER metal4 ;
  RECT 3612.860 1356.100 3613.980 1359.340 ;
  LAYER metal3 ;
  RECT 3612.860 1356.100 3613.980 1359.340 ;
  LAYER metal2 ;
  RECT 3612.860 1356.100 3613.980 1359.340 ;
  LAYER metal1 ;
  RECT 3612.860 1356.100 3613.980 1359.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1348.260 3613.980 1351.500 ;
  LAYER metal4 ;
  RECT 3612.860 1348.260 3613.980 1351.500 ;
  LAYER metal3 ;
  RECT 3612.860 1348.260 3613.980 1351.500 ;
  LAYER metal2 ;
  RECT 3612.860 1348.260 3613.980 1351.500 ;
  LAYER metal1 ;
  RECT 3612.860 1348.260 3613.980 1351.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1340.420 3613.980 1343.660 ;
  LAYER metal4 ;
  RECT 3612.860 1340.420 3613.980 1343.660 ;
  LAYER metal3 ;
  RECT 3612.860 1340.420 3613.980 1343.660 ;
  LAYER metal2 ;
  RECT 3612.860 1340.420 3613.980 1343.660 ;
  LAYER metal1 ;
  RECT 3612.860 1340.420 3613.980 1343.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1301.220 3613.980 1304.460 ;
  LAYER metal4 ;
  RECT 3612.860 1301.220 3613.980 1304.460 ;
  LAYER metal3 ;
  RECT 3612.860 1301.220 3613.980 1304.460 ;
  LAYER metal2 ;
  RECT 3612.860 1301.220 3613.980 1304.460 ;
  LAYER metal1 ;
  RECT 3612.860 1301.220 3613.980 1304.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1293.380 3613.980 1296.620 ;
  LAYER metal4 ;
  RECT 3612.860 1293.380 3613.980 1296.620 ;
  LAYER metal3 ;
  RECT 3612.860 1293.380 3613.980 1296.620 ;
  LAYER metal2 ;
  RECT 3612.860 1293.380 3613.980 1296.620 ;
  LAYER metal1 ;
  RECT 3612.860 1293.380 3613.980 1296.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1285.540 3613.980 1288.780 ;
  LAYER metal4 ;
  RECT 3612.860 1285.540 3613.980 1288.780 ;
  LAYER metal3 ;
  RECT 3612.860 1285.540 3613.980 1288.780 ;
  LAYER metal2 ;
  RECT 3612.860 1285.540 3613.980 1288.780 ;
  LAYER metal1 ;
  RECT 3612.860 1285.540 3613.980 1288.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1277.700 3613.980 1280.940 ;
  LAYER metal4 ;
  RECT 3612.860 1277.700 3613.980 1280.940 ;
  LAYER metal3 ;
  RECT 3612.860 1277.700 3613.980 1280.940 ;
  LAYER metal2 ;
  RECT 3612.860 1277.700 3613.980 1280.940 ;
  LAYER metal1 ;
  RECT 3612.860 1277.700 3613.980 1280.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1269.860 3613.980 1273.100 ;
  LAYER metal4 ;
  RECT 3612.860 1269.860 3613.980 1273.100 ;
  LAYER metal3 ;
  RECT 3612.860 1269.860 3613.980 1273.100 ;
  LAYER metal2 ;
  RECT 3612.860 1269.860 3613.980 1273.100 ;
  LAYER metal1 ;
  RECT 3612.860 1269.860 3613.980 1273.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1262.020 3613.980 1265.260 ;
  LAYER metal4 ;
  RECT 3612.860 1262.020 3613.980 1265.260 ;
  LAYER metal3 ;
  RECT 3612.860 1262.020 3613.980 1265.260 ;
  LAYER metal2 ;
  RECT 3612.860 1262.020 3613.980 1265.260 ;
  LAYER metal1 ;
  RECT 3612.860 1262.020 3613.980 1265.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1222.820 3613.980 1226.060 ;
  LAYER metal4 ;
  RECT 3612.860 1222.820 3613.980 1226.060 ;
  LAYER metal3 ;
  RECT 3612.860 1222.820 3613.980 1226.060 ;
  LAYER metal2 ;
  RECT 3612.860 1222.820 3613.980 1226.060 ;
  LAYER metal1 ;
  RECT 3612.860 1222.820 3613.980 1226.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1214.980 3613.980 1218.220 ;
  LAYER metal4 ;
  RECT 3612.860 1214.980 3613.980 1218.220 ;
  LAYER metal3 ;
  RECT 3612.860 1214.980 3613.980 1218.220 ;
  LAYER metal2 ;
  RECT 3612.860 1214.980 3613.980 1218.220 ;
  LAYER metal1 ;
  RECT 3612.860 1214.980 3613.980 1218.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1207.140 3613.980 1210.380 ;
  LAYER metal4 ;
  RECT 3612.860 1207.140 3613.980 1210.380 ;
  LAYER metal3 ;
  RECT 3612.860 1207.140 3613.980 1210.380 ;
  LAYER metal2 ;
  RECT 3612.860 1207.140 3613.980 1210.380 ;
  LAYER metal1 ;
  RECT 3612.860 1207.140 3613.980 1210.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1199.300 3613.980 1202.540 ;
  LAYER metal4 ;
  RECT 3612.860 1199.300 3613.980 1202.540 ;
  LAYER metal3 ;
  RECT 3612.860 1199.300 3613.980 1202.540 ;
  LAYER metal2 ;
  RECT 3612.860 1199.300 3613.980 1202.540 ;
  LAYER metal1 ;
  RECT 3612.860 1199.300 3613.980 1202.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1191.460 3613.980 1194.700 ;
  LAYER metal4 ;
  RECT 3612.860 1191.460 3613.980 1194.700 ;
  LAYER metal3 ;
  RECT 3612.860 1191.460 3613.980 1194.700 ;
  LAYER metal2 ;
  RECT 3612.860 1191.460 3613.980 1194.700 ;
  LAYER metal1 ;
  RECT 3612.860 1191.460 3613.980 1194.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1183.620 3613.980 1186.860 ;
  LAYER metal4 ;
  RECT 3612.860 1183.620 3613.980 1186.860 ;
  LAYER metal3 ;
  RECT 3612.860 1183.620 3613.980 1186.860 ;
  LAYER metal2 ;
  RECT 3612.860 1183.620 3613.980 1186.860 ;
  LAYER metal1 ;
  RECT 3612.860 1183.620 3613.980 1186.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1144.420 3613.980 1147.660 ;
  LAYER metal4 ;
  RECT 3612.860 1144.420 3613.980 1147.660 ;
  LAYER metal3 ;
  RECT 3612.860 1144.420 3613.980 1147.660 ;
  LAYER metal2 ;
  RECT 3612.860 1144.420 3613.980 1147.660 ;
  LAYER metal1 ;
  RECT 3612.860 1144.420 3613.980 1147.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1136.580 3613.980 1139.820 ;
  LAYER metal4 ;
  RECT 3612.860 1136.580 3613.980 1139.820 ;
  LAYER metal3 ;
  RECT 3612.860 1136.580 3613.980 1139.820 ;
  LAYER metal2 ;
  RECT 3612.860 1136.580 3613.980 1139.820 ;
  LAYER metal1 ;
  RECT 3612.860 1136.580 3613.980 1139.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1128.740 3613.980 1131.980 ;
  LAYER metal4 ;
  RECT 3612.860 1128.740 3613.980 1131.980 ;
  LAYER metal3 ;
  RECT 3612.860 1128.740 3613.980 1131.980 ;
  LAYER metal2 ;
  RECT 3612.860 1128.740 3613.980 1131.980 ;
  LAYER metal1 ;
  RECT 3612.860 1128.740 3613.980 1131.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1120.900 3613.980 1124.140 ;
  LAYER metal4 ;
  RECT 3612.860 1120.900 3613.980 1124.140 ;
  LAYER metal3 ;
  RECT 3612.860 1120.900 3613.980 1124.140 ;
  LAYER metal2 ;
  RECT 3612.860 1120.900 3613.980 1124.140 ;
  LAYER metal1 ;
  RECT 3612.860 1120.900 3613.980 1124.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1113.060 3613.980 1116.300 ;
  LAYER metal4 ;
  RECT 3612.860 1113.060 3613.980 1116.300 ;
  LAYER metal3 ;
  RECT 3612.860 1113.060 3613.980 1116.300 ;
  LAYER metal2 ;
  RECT 3612.860 1113.060 3613.980 1116.300 ;
  LAYER metal1 ;
  RECT 3612.860 1113.060 3613.980 1116.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1105.220 3613.980 1108.460 ;
  LAYER metal4 ;
  RECT 3612.860 1105.220 3613.980 1108.460 ;
  LAYER metal3 ;
  RECT 3612.860 1105.220 3613.980 1108.460 ;
  LAYER metal2 ;
  RECT 3612.860 1105.220 3613.980 1108.460 ;
  LAYER metal1 ;
  RECT 3612.860 1105.220 3613.980 1108.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1066.020 3613.980 1069.260 ;
  LAYER metal4 ;
  RECT 3612.860 1066.020 3613.980 1069.260 ;
  LAYER metal3 ;
  RECT 3612.860 1066.020 3613.980 1069.260 ;
  LAYER metal2 ;
  RECT 3612.860 1066.020 3613.980 1069.260 ;
  LAYER metal1 ;
  RECT 3612.860 1066.020 3613.980 1069.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1058.180 3613.980 1061.420 ;
  LAYER metal4 ;
  RECT 3612.860 1058.180 3613.980 1061.420 ;
  LAYER metal3 ;
  RECT 3612.860 1058.180 3613.980 1061.420 ;
  LAYER metal2 ;
  RECT 3612.860 1058.180 3613.980 1061.420 ;
  LAYER metal1 ;
  RECT 3612.860 1058.180 3613.980 1061.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1050.340 3613.980 1053.580 ;
  LAYER metal4 ;
  RECT 3612.860 1050.340 3613.980 1053.580 ;
  LAYER metal3 ;
  RECT 3612.860 1050.340 3613.980 1053.580 ;
  LAYER metal2 ;
  RECT 3612.860 1050.340 3613.980 1053.580 ;
  LAYER metal1 ;
  RECT 3612.860 1050.340 3613.980 1053.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1042.500 3613.980 1045.740 ;
  LAYER metal4 ;
  RECT 3612.860 1042.500 3613.980 1045.740 ;
  LAYER metal3 ;
  RECT 3612.860 1042.500 3613.980 1045.740 ;
  LAYER metal2 ;
  RECT 3612.860 1042.500 3613.980 1045.740 ;
  LAYER metal1 ;
  RECT 3612.860 1042.500 3613.980 1045.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1034.660 3613.980 1037.900 ;
  LAYER metal4 ;
  RECT 3612.860 1034.660 3613.980 1037.900 ;
  LAYER metal3 ;
  RECT 3612.860 1034.660 3613.980 1037.900 ;
  LAYER metal2 ;
  RECT 3612.860 1034.660 3613.980 1037.900 ;
  LAYER metal1 ;
  RECT 3612.860 1034.660 3613.980 1037.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 1026.820 3613.980 1030.060 ;
  LAYER metal4 ;
  RECT 3612.860 1026.820 3613.980 1030.060 ;
  LAYER metal3 ;
  RECT 3612.860 1026.820 3613.980 1030.060 ;
  LAYER metal2 ;
  RECT 3612.860 1026.820 3613.980 1030.060 ;
  LAYER metal1 ;
  RECT 3612.860 1026.820 3613.980 1030.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 987.620 3613.980 990.860 ;
  LAYER metal4 ;
  RECT 3612.860 987.620 3613.980 990.860 ;
  LAYER metal3 ;
  RECT 3612.860 987.620 3613.980 990.860 ;
  LAYER metal2 ;
  RECT 3612.860 987.620 3613.980 990.860 ;
  LAYER metal1 ;
  RECT 3612.860 987.620 3613.980 990.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 979.780 3613.980 983.020 ;
  LAYER metal4 ;
  RECT 3612.860 979.780 3613.980 983.020 ;
  LAYER metal3 ;
  RECT 3612.860 979.780 3613.980 983.020 ;
  LAYER metal2 ;
  RECT 3612.860 979.780 3613.980 983.020 ;
  LAYER metal1 ;
  RECT 3612.860 979.780 3613.980 983.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 971.940 3613.980 975.180 ;
  LAYER metal4 ;
  RECT 3612.860 971.940 3613.980 975.180 ;
  LAYER metal3 ;
  RECT 3612.860 971.940 3613.980 975.180 ;
  LAYER metal2 ;
  RECT 3612.860 971.940 3613.980 975.180 ;
  LAYER metal1 ;
  RECT 3612.860 971.940 3613.980 975.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 964.100 3613.980 967.340 ;
  LAYER metal4 ;
  RECT 3612.860 964.100 3613.980 967.340 ;
  LAYER metal3 ;
  RECT 3612.860 964.100 3613.980 967.340 ;
  LAYER metal2 ;
  RECT 3612.860 964.100 3613.980 967.340 ;
  LAYER metal1 ;
  RECT 3612.860 964.100 3613.980 967.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 956.260 3613.980 959.500 ;
  LAYER metal4 ;
  RECT 3612.860 956.260 3613.980 959.500 ;
  LAYER metal3 ;
  RECT 3612.860 956.260 3613.980 959.500 ;
  LAYER metal2 ;
  RECT 3612.860 956.260 3613.980 959.500 ;
  LAYER metal1 ;
  RECT 3612.860 956.260 3613.980 959.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 948.420 3613.980 951.660 ;
  LAYER metal4 ;
  RECT 3612.860 948.420 3613.980 951.660 ;
  LAYER metal3 ;
  RECT 3612.860 948.420 3613.980 951.660 ;
  LAYER metal2 ;
  RECT 3612.860 948.420 3613.980 951.660 ;
  LAYER metal1 ;
  RECT 3612.860 948.420 3613.980 951.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 909.220 3613.980 912.460 ;
  LAYER metal4 ;
  RECT 3612.860 909.220 3613.980 912.460 ;
  LAYER metal3 ;
  RECT 3612.860 909.220 3613.980 912.460 ;
  LAYER metal2 ;
  RECT 3612.860 909.220 3613.980 912.460 ;
  LAYER metal1 ;
  RECT 3612.860 909.220 3613.980 912.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 901.380 3613.980 904.620 ;
  LAYER metal4 ;
  RECT 3612.860 901.380 3613.980 904.620 ;
  LAYER metal3 ;
  RECT 3612.860 901.380 3613.980 904.620 ;
  LAYER metal2 ;
  RECT 3612.860 901.380 3613.980 904.620 ;
  LAYER metal1 ;
  RECT 3612.860 901.380 3613.980 904.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 893.540 3613.980 896.780 ;
  LAYER metal4 ;
  RECT 3612.860 893.540 3613.980 896.780 ;
  LAYER metal3 ;
  RECT 3612.860 893.540 3613.980 896.780 ;
  LAYER metal2 ;
  RECT 3612.860 893.540 3613.980 896.780 ;
  LAYER metal1 ;
  RECT 3612.860 893.540 3613.980 896.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 885.700 3613.980 888.940 ;
  LAYER metal4 ;
  RECT 3612.860 885.700 3613.980 888.940 ;
  LAYER metal3 ;
  RECT 3612.860 885.700 3613.980 888.940 ;
  LAYER metal2 ;
  RECT 3612.860 885.700 3613.980 888.940 ;
  LAYER metal1 ;
  RECT 3612.860 885.700 3613.980 888.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 877.860 3613.980 881.100 ;
  LAYER metal4 ;
  RECT 3612.860 877.860 3613.980 881.100 ;
  LAYER metal3 ;
  RECT 3612.860 877.860 3613.980 881.100 ;
  LAYER metal2 ;
  RECT 3612.860 877.860 3613.980 881.100 ;
  LAYER metal1 ;
  RECT 3612.860 877.860 3613.980 881.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 870.020 3613.980 873.260 ;
  LAYER metal4 ;
  RECT 3612.860 870.020 3613.980 873.260 ;
  LAYER metal3 ;
  RECT 3612.860 870.020 3613.980 873.260 ;
  LAYER metal2 ;
  RECT 3612.860 870.020 3613.980 873.260 ;
  LAYER metal1 ;
  RECT 3612.860 870.020 3613.980 873.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 830.820 3613.980 834.060 ;
  LAYER metal4 ;
  RECT 3612.860 830.820 3613.980 834.060 ;
  LAYER metal3 ;
  RECT 3612.860 830.820 3613.980 834.060 ;
  LAYER metal2 ;
  RECT 3612.860 830.820 3613.980 834.060 ;
  LAYER metal1 ;
  RECT 3612.860 830.820 3613.980 834.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 822.980 3613.980 826.220 ;
  LAYER metal4 ;
  RECT 3612.860 822.980 3613.980 826.220 ;
  LAYER metal3 ;
  RECT 3612.860 822.980 3613.980 826.220 ;
  LAYER metal2 ;
  RECT 3612.860 822.980 3613.980 826.220 ;
  LAYER metal1 ;
  RECT 3612.860 822.980 3613.980 826.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 815.140 3613.980 818.380 ;
  LAYER metal4 ;
  RECT 3612.860 815.140 3613.980 818.380 ;
  LAYER metal3 ;
  RECT 3612.860 815.140 3613.980 818.380 ;
  LAYER metal2 ;
  RECT 3612.860 815.140 3613.980 818.380 ;
  LAYER metal1 ;
  RECT 3612.860 815.140 3613.980 818.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 807.300 3613.980 810.540 ;
  LAYER metal4 ;
  RECT 3612.860 807.300 3613.980 810.540 ;
  LAYER metal3 ;
  RECT 3612.860 807.300 3613.980 810.540 ;
  LAYER metal2 ;
  RECT 3612.860 807.300 3613.980 810.540 ;
  LAYER metal1 ;
  RECT 3612.860 807.300 3613.980 810.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 799.460 3613.980 802.700 ;
  LAYER metal4 ;
  RECT 3612.860 799.460 3613.980 802.700 ;
  LAYER metal3 ;
  RECT 3612.860 799.460 3613.980 802.700 ;
  LAYER metal2 ;
  RECT 3612.860 799.460 3613.980 802.700 ;
  LAYER metal1 ;
  RECT 3612.860 799.460 3613.980 802.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 791.620 3613.980 794.860 ;
  LAYER metal4 ;
  RECT 3612.860 791.620 3613.980 794.860 ;
  LAYER metal3 ;
  RECT 3612.860 791.620 3613.980 794.860 ;
  LAYER metal2 ;
  RECT 3612.860 791.620 3613.980 794.860 ;
  LAYER metal1 ;
  RECT 3612.860 791.620 3613.980 794.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 752.420 3613.980 755.660 ;
  LAYER metal4 ;
  RECT 3612.860 752.420 3613.980 755.660 ;
  LAYER metal3 ;
  RECT 3612.860 752.420 3613.980 755.660 ;
  LAYER metal2 ;
  RECT 3612.860 752.420 3613.980 755.660 ;
  LAYER metal1 ;
  RECT 3612.860 752.420 3613.980 755.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 744.580 3613.980 747.820 ;
  LAYER metal4 ;
  RECT 3612.860 744.580 3613.980 747.820 ;
  LAYER metal3 ;
  RECT 3612.860 744.580 3613.980 747.820 ;
  LAYER metal2 ;
  RECT 3612.860 744.580 3613.980 747.820 ;
  LAYER metal1 ;
  RECT 3612.860 744.580 3613.980 747.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 736.740 3613.980 739.980 ;
  LAYER metal4 ;
  RECT 3612.860 736.740 3613.980 739.980 ;
  LAYER metal3 ;
  RECT 3612.860 736.740 3613.980 739.980 ;
  LAYER metal2 ;
  RECT 3612.860 736.740 3613.980 739.980 ;
  LAYER metal1 ;
  RECT 3612.860 736.740 3613.980 739.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 728.900 3613.980 732.140 ;
  LAYER metal4 ;
  RECT 3612.860 728.900 3613.980 732.140 ;
  LAYER metal3 ;
  RECT 3612.860 728.900 3613.980 732.140 ;
  LAYER metal2 ;
  RECT 3612.860 728.900 3613.980 732.140 ;
  LAYER metal1 ;
  RECT 3612.860 728.900 3613.980 732.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 721.060 3613.980 724.300 ;
  LAYER metal4 ;
  RECT 3612.860 721.060 3613.980 724.300 ;
  LAYER metal3 ;
  RECT 3612.860 721.060 3613.980 724.300 ;
  LAYER metal2 ;
  RECT 3612.860 721.060 3613.980 724.300 ;
  LAYER metal1 ;
  RECT 3612.860 721.060 3613.980 724.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 713.220 3613.980 716.460 ;
  LAYER metal4 ;
  RECT 3612.860 713.220 3613.980 716.460 ;
  LAYER metal3 ;
  RECT 3612.860 713.220 3613.980 716.460 ;
  LAYER metal2 ;
  RECT 3612.860 713.220 3613.980 716.460 ;
  LAYER metal1 ;
  RECT 3612.860 713.220 3613.980 716.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 674.020 3613.980 677.260 ;
  LAYER metal4 ;
  RECT 3612.860 674.020 3613.980 677.260 ;
  LAYER metal3 ;
  RECT 3612.860 674.020 3613.980 677.260 ;
  LAYER metal2 ;
  RECT 3612.860 674.020 3613.980 677.260 ;
  LAYER metal1 ;
  RECT 3612.860 674.020 3613.980 677.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 666.180 3613.980 669.420 ;
  LAYER metal4 ;
  RECT 3612.860 666.180 3613.980 669.420 ;
  LAYER metal3 ;
  RECT 3612.860 666.180 3613.980 669.420 ;
  LAYER metal2 ;
  RECT 3612.860 666.180 3613.980 669.420 ;
  LAYER metal1 ;
  RECT 3612.860 666.180 3613.980 669.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 658.340 3613.980 661.580 ;
  LAYER metal4 ;
  RECT 3612.860 658.340 3613.980 661.580 ;
  LAYER metal3 ;
  RECT 3612.860 658.340 3613.980 661.580 ;
  LAYER metal2 ;
  RECT 3612.860 658.340 3613.980 661.580 ;
  LAYER metal1 ;
  RECT 3612.860 658.340 3613.980 661.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 650.500 3613.980 653.740 ;
  LAYER metal4 ;
  RECT 3612.860 650.500 3613.980 653.740 ;
  LAYER metal3 ;
  RECT 3612.860 650.500 3613.980 653.740 ;
  LAYER metal2 ;
  RECT 3612.860 650.500 3613.980 653.740 ;
  LAYER metal1 ;
  RECT 3612.860 650.500 3613.980 653.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 642.660 3613.980 645.900 ;
  LAYER metal4 ;
  RECT 3612.860 642.660 3613.980 645.900 ;
  LAYER metal3 ;
  RECT 3612.860 642.660 3613.980 645.900 ;
  LAYER metal2 ;
  RECT 3612.860 642.660 3613.980 645.900 ;
  LAYER metal1 ;
  RECT 3612.860 642.660 3613.980 645.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 634.820 3613.980 638.060 ;
  LAYER metal4 ;
  RECT 3612.860 634.820 3613.980 638.060 ;
  LAYER metal3 ;
  RECT 3612.860 634.820 3613.980 638.060 ;
  LAYER metal2 ;
  RECT 3612.860 634.820 3613.980 638.060 ;
  LAYER metal1 ;
  RECT 3612.860 634.820 3613.980 638.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 595.620 3613.980 598.860 ;
  LAYER metal4 ;
  RECT 3612.860 595.620 3613.980 598.860 ;
  LAYER metal3 ;
  RECT 3612.860 595.620 3613.980 598.860 ;
  LAYER metal2 ;
  RECT 3612.860 595.620 3613.980 598.860 ;
  LAYER metal1 ;
  RECT 3612.860 595.620 3613.980 598.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 587.780 3613.980 591.020 ;
  LAYER metal4 ;
  RECT 3612.860 587.780 3613.980 591.020 ;
  LAYER metal3 ;
  RECT 3612.860 587.780 3613.980 591.020 ;
  LAYER metal2 ;
  RECT 3612.860 587.780 3613.980 591.020 ;
  LAYER metal1 ;
  RECT 3612.860 587.780 3613.980 591.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 579.940 3613.980 583.180 ;
  LAYER metal4 ;
  RECT 3612.860 579.940 3613.980 583.180 ;
  LAYER metal3 ;
  RECT 3612.860 579.940 3613.980 583.180 ;
  LAYER metal2 ;
  RECT 3612.860 579.940 3613.980 583.180 ;
  LAYER metal1 ;
  RECT 3612.860 579.940 3613.980 583.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 572.100 3613.980 575.340 ;
  LAYER metal4 ;
  RECT 3612.860 572.100 3613.980 575.340 ;
  LAYER metal3 ;
  RECT 3612.860 572.100 3613.980 575.340 ;
  LAYER metal2 ;
  RECT 3612.860 572.100 3613.980 575.340 ;
  LAYER metal1 ;
  RECT 3612.860 572.100 3613.980 575.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 564.260 3613.980 567.500 ;
  LAYER metal4 ;
  RECT 3612.860 564.260 3613.980 567.500 ;
  LAYER metal3 ;
  RECT 3612.860 564.260 3613.980 567.500 ;
  LAYER metal2 ;
  RECT 3612.860 564.260 3613.980 567.500 ;
  LAYER metal1 ;
  RECT 3612.860 564.260 3613.980 567.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 556.420 3613.980 559.660 ;
  LAYER metal4 ;
  RECT 3612.860 556.420 3613.980 559.660 ;
  LAYER metal3 ;
  RECT 3612.860 556.420 3613.980 559.660 ;
  LAYER metal2 ;
  RECT 3612.860 556.420 3613.980 559.660 ;
  LAYER metal1 ;
  RECT 3612.860 556.420 3613.980 559.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 517.220 3613.980 520.460 ;
  LAYER metal4 ;
  RECT 3612.860 517.220 3613.980 520.460 ;
  LAYER metal3 ;
  RECT 3612.860 517.220 3613.980 520.460 ;
  LAYER metal2 ;
  RECT 3612.860 517.220 3613.980 520.460 ;
  LAYER metal1 ;
  RECT 3612.860 517.220 3613.980 520.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 509.380 3613.980 512.620 ;
  LAYER metal4 ;
  RECT 3612.860 509.380 3613.980 512.620 ;
  LAYER metal3 ;
  RECT 3612.860 509.380 3613.980 512.620 ;
  LAYER metal2 ;
  RECT 3612.860 509.380 3613.980 512.620 ;
  LAYER metal1 ;
  RECT 3612.860 509.380 3613.980 512.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 501.540 3613.980 504.780 ;
  LAYER metal4 ;
  RECT 3612.860 501.540 3613.980 504.780 ;
  LAYER metal3 ;
  RECT 3612.860 501.540 3613.980 504.780 ;
  LAYER metal2 ;
  RECT 3612.860 501.540 3613.980 504.780 ;
  LAYER metal1 ;
  RECT 3612.860 501.540 3613.980 504.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 493.700 3613.980 496.940 ;
  LAYER metal4 ;
  RECT 3612.860 493.700 3613.980 496.940 ;
  LAYER metal3 ;
  RECT 3612.860 493.700 3613.980 496.940 ;
  LAYER metal2 ;
  RECT 3612.860 493.700 3613.980 496.940 ;
  LAYER metal1 ;
  RECT 3612.860 493.700 3613.980 496.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 485.860 3613.980 489.100 ;
  LAYER metal4 ;
  RECT 3612.860 485.860 3613.980 489.100 ;
  LAYER metal3 ;
  RECT 3612.860 485.860 3613.980 489.100 ;
  LAYER metal2 ;
  RECT 3612.860 485.860 3613.980 489.100 ;
  LAYER metal1 ;
  RECT 3612.860 485.860 3613.980 489.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 478.020 3613.980 481.260 ;
  LAYER metal4 ;
  RECT 3612.860 478.020 3613.980 481.260 ;
  LAYER metal3 ;
  RECT 3612.860 478.020 3613.980 481.260 ;
  LAYER metal2 ;
  RECT 3612.860 478.020 3613.980 481.260 ;
  LAYER metal1 ;
  RECT 3612.860 478.020 3613.980 481.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 438.820 3613.980 442.060 ;
  LAYER metal4 ;
  RECT 3612.860 438.820 3613.980 442.060 ;
  LAYER metal3 ;
  RECT 3612.860 438.820 3613.980 442.060 ;
  LAYER metal2 ;
  RECT 3612.860 438.820 3613.980 442.060 ;
  LAYER metal1 ;
  RECT 3612.860 438.820 3613.980 442.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 430.980 3613.980 434.220 ;
  LAYER metal4 ;
  RECT 3612.860 430.980 3613.980 434.220 ;
  LAYER metal3 ;
  RECT 3612.860 430.980 3613.980 434.220 ;
  LAYER metal2 ;
  RECT 3612.860 430.980 3613.980 434.220 ;
  LAYER metal1 ;
  RECT 3612.860 430.980 3613.980 434.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 423.140 3613.980 426.380 ;
  LAYER metal4 ;
  RECT 3612.860 423.140 3613.980 426.380 ;
  LAYER metal3 ;
  RECT 3612.860 423.140 3613.980 426.380 ;
  LAYER metal2 ;
  RECT 3612.860 423.140 3613.980 426.380 ;
  LAYER metal1 ;
  RECT 3612.860 423.140 3613.980 426.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 415.300 3613.980 418.540 ;
  LAYER metal4 ;
  RECT 3612.860 415.300 3613.980 418.540 ;
  LAYER metal3 ;
  RECT 3612.860 415.300 3613.980 418.540 ;
  LAYER metal2 ;
  RECT 3612.860 415.300 3613.980 418.540 ;
  LAYER metal1 ;
  RECT 3612.860 415.300 3613.980 418.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 407.460 3613.980 410.700 ;
  LAYER metal4 ;
  RECT 3612.860 407.460 3613.980 410.700 ;
  LAYER metal3 ;
  RECT 3612.860 407.460 3613.980 410.700 ;
  LAYER metal2 ;
  RECT 3612.860 407.460 3613.980 410.700 ;
  LAYER metal1 ;
  RECT 3612.860 407.460 3613.980 410.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 399.620 3613.980 402.860 ;
  LAYER metal4 ;
  RECT 3612.860 399.620 3613.980 402.860 ;
  LAYER metal3 ;
  RECT 3612.860 399.620 3613.980 402.860 ;
  LAYER metal2 ;
  RECT 3612.860 399.620 3613.980 402.860 ;
  LAYER metal1 ;
  RECT 3612.860 399.620 3613.980 402.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 360.420 3613.980 363.660 ;
  LAYER metal4 ;
  RECT 3612.860 360.420 3613.980 363.660 ;
  LAYER metal3 ;
  RECT 3612.860 360.420 3613.980 363.660 ;
  LAYER metal2 ;
  RECT 3612.860 360.420 3613.980 363.660 ;
  LAYER metal1 ;
  RECT 3612.860 360.420 3613.980 363.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 352.580 3613.980 355.820 ;
  LAYER metal4 ;
  RECT 3612.860 352.580 3613.980 355.820 ;
  LAYER metal3 ;
  RECT 3612.860 352.580 3613.980 355.820 ;
  LAYER metal2 ;
  RECT 3612.860 352.580 3613.980 355.820 ;
  LAYER metal1 ;
  RECT 3612.860 352.580 3613.980 355.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 344.740 3613.980 347.980 ;
  LAYER metal4 ;
  RECT 3612.860 344.740 3613.980 347.980 ;
  LAYER metal3 ;
  RECT 3612.860 344.740 3613.980 347.980 ;
  LAYER metal2 ;
  RECT 3612.860 344.740 3613.980 347.980 ;
  LAYER metal1 ;
  RECT 3612.860 344.740 3613.980 347.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 336.900 3613.980 340.140 ;
  LAYER metal4 ;
  RECT 3612.860 336.900 3613.980 340.140 ;
  LAYER metal3 ;
  RECT 3612.860 336.900 3613.980 340.140 ;
  LAYER metal2 ;
  RECT 3612.860 336.900 3613.980 340.140 ;
  LAYER metal1 ;
  RECT 3612.860 336.900 3613.980 340.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 329.060 3613.980 332.300 ;
  LAYER metal4 ;
  RECT 3612.860 329.060 3613.980 332.300 ;
  LAYER metal3 ;
  RECT 3612.860 329.060 3613.980 332.300 ;
  LAYER metal2 ;
  RECT 3612.860 329.060 3613.980 332.300 ;
  LAYER metal1 ;
  RECT 3612.860 329.060 3613.980 332.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 321.220 3613.980 324.460 ;
  LAYER metal4 ;
  RECT 3612.860 321.220 3613.980 324.460 ;
  LAYER metal3 ;
  RECT 3612.860 321.220 3613.980 324.460 ;
  LAYER metal2 ;
  RECT 3612.860 321.220 3613.980 324.460 ;
  LAYER metal1 ;
  RECT 3612.860 321.220 3613.980 324.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 282.020 3613.980 285.260 ;
  LAYER metal4 ;
  RECT 3612.860 282.020 3613.980 285.260 ;
  LAYER metal3 ;
  RECT 3612.860 282.020 3613.980 285.260 ;
  LAYER metal2 ;
  RECT 3612.860 282.020 3613.980 285.260 ;
  LAYER metal1 ;
  RECT 3612.860 282.020 3613.980 285.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 274.180 3613.980 277.420 ;
  LAYER metal4 ;
  RECT 3612.860 274.180 3613.980 277.420 ;
  LAYER metal3 ;
  RECT 3612.860 274.180 3613.980 277.420 ;
  LAYER metal2 ;
  RECT 3612.860 274.180 3613.980 277.420 ;
  LAYER metal1 ;
  RECT 3612.860 274.180 3613.980 277.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 266.340 3613.980 269.580 ;
  LAYER metal4 ;
  RECT 3612.860 266.340 3613.980 269.580 ;
  LAYER metal3 ;
  RECT 3612.860 266.340 3613.980 269.580 ;
  LAYER metal2 ;
  RECT 3612.860 266.340 3613.980 269.580 ;
  LAYER metal1 ;
  RECT 3612.860 266.340 3613.980 269.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 258.500 3613.980 261.740 ;
  LAYER metal4 ;
  RECT 3612.860 258.500 3613.980 261.740 ;
  LAYER metal3 ;
  RECT 3612.860 258.500 3613.980 261.740 ;
  LAYER metal2 ;
  RECT 3612.860 258.500 3613.980 261.740 ;
  LAYER metal1 ;
  RECT 3612.860 258.500 3613.980 261.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 250.660 3613.980 253.900 ;
  LAYER metal4 ;
  RECT 3612.860 250.660 3613.980 253.900 ;
  LAYER metal3 ;
  RECT 3612.860 250.660 3613.980 253.900 ;
  LAYER metal2 ;
  RECT 3612.860 250.660 3613.980 253.900 ;
  LAYER metal1 ;
  RECT 3612.860 250.660 3613.980 253.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 242.820 3613.980 246.060 ;
  LAYER metal4 ;
  RECT 3612.860 242.820 3613.980 246.060 ;
  LAYER metal3 ;
  RECT 3612.860 242.820 3613.980 246.060 ;
  LAYER metal2 ;
  RECT 3612.860 242.820 3613.980 246.060 ;
  LAYER metal1 ;
  RECT 3612.860 242.820 3613.980 246.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 203.620 3613.980 206.860 ;
  LAYER metal4 ;
  RECT 3612.860 203.620 3613.980 206.860 ;
  LAYER metal3 ;
  RECT 3612.860 203.620 3613.980 206.860 ;
  LAYER metal2 ;
  RECT 3612.860 203.620 3613.980 206.860 ;
  LAYER metal1 ;
  RECT 3612.860 203.620 3613.980 206.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 195.780 3613.980 199.020 ;
  LAYER metal4 ;
  RECT 3612.860 195.780 3613.980 199.020 ;
  LAYER metal3 ;
  RECT 3612.860 195.780 3613.980 199.020 ;
  LAYER metal2 ;
  RECT 3612.860 195.780 3613.980 199.020 ;
  LAYER metal1 ;
  RECT 3612.860 195.780 3613.980 199.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 187.940 3613.980 191.180 ;
  LAYER metal4 ;
  RECT 3612.860 187.940 3613.980 191.180 ;
  LAYER metal3 ;
  RECT 3612.860 187.940 3613.980 191.180 ;
  LAYER metal2 ;
  RECT 3612.860 187.940 3613.980 191.180 ;
  LAYER metal1 ;
  RECT 3612.860 187.940 3613.980 191.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 180.100 3613.980 183.340 ;
  LAYER metal4 ;
  RECT 3612.860 180.100 3613.980 183.340 ;
  LAYER metal3 ;
  RECT 3612.860 180.100 3613.980 183.340 ;
  LAYER metal2 ;
  RECT 3612.860 180.100 3613.980 183.340 ;
  LAYER metal1 ;
  RECT 3612.860 180.100 3613.980 183.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 172.260 3613.980 175.500 ;
  LAYER metal4 ;
  RECT 3612.860 172.260 3613.980 175.500 ;
  LAYER metal3 ;
  RECT 3612.860 172.260 3613.980 175.500 ;
  LAYER metal2 ;
  RECT 3612.860 172.260 3613.980 175.500 ;
  LAYER metal1 ;
  RECT 3612.860 172.260 3613.980 175.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 164.420 3613.980 167.660 ;
  LAYER metal4 ;
  RECT 3612.860 164.420 3613.980 167.660 ;
  LAYER metal3 ;
  RECT 3612.860 164.420 3613.980 167.660 ;
  LAYER metal2 ;
  RECT 3612.860 164.420 3613.980 167.660 ;
  LAYER metal1 ;
  RECT 3612.860 164.420 3613.980 167.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 125.220 3613.980 128.460 ;
  LAYER metal4 ;
  RECT 3612.860 125.220 3613.980 128.460 ;
  LAYER metal3 ;
  RECT 3612.860 125.220 3613.980 128.460 ;
  LAYER metal2 ;
  RECT 3612.860 125.220 3613.980 128.460 ;
  LAYER metal1 ;
  RECT 3612.860 125.220 3613.980 128.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 117.380 3613.980 120.620 ;
  LAYER metal4 ;
  RECT 3612.860 117.380 3613.980 120.620 ;
  LAYER metal3 ;
  RECT 3612.860 117.380 3613.980 120.620 ;
  LAYER metal2 ;
  RECT 3612.860 117.380 3613.980 120.620 ;
  LAYER metal1 ;
  RECT 3612.860 117.380 3613.980 120.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 109.540 3613.980 112.780 ;
  LAYER metal4 ;
  RECT 3612.860 109.540 3613.980 112.780 ;
  LAYER metal3 ;
  RECT 3612.860 109.540 3613.980 112.780 ;
  LAYER metal2 ;
  RECT 3612.860 109.540 3613.980 112.780 ;
  LAYER metal1 ;
  RECT 3612.860 109.540 3613.980 112.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 101.700 3613.980 104.940 ;
  LAYER metal4 ;
  RECT 3612.860 101.700 3613.980 104.940 ;
  LAYER metal3 ;
  RECT 3612.860 101.700 3613.980 104.940 ;
  LAYER metal2 ;
  RECT 3612.860 101.700 3613.980 104.940 ;
  LAYER metal1 ;
  RECT 3612.860 101.700 3613.980 104.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 93.860 3613.980 97.100 ;
  LAYER metal4 ;
  RECT 3612.860 93.860 3613.980 97.100 ;
  LAYER metal3 ;
  RECT 3612.860 93.860 3613.980 97.100 ;
  LAYER metal2 ;
  RECT 3612.860 93.860 3613.980 97.100 ;
  LAYER metal1 ;
  RECT 3612.860 93.860 3613.980 97.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 86.020 3613.980 89.260 ;
  LAYER metal4 ;
  RECT 3612.860 86.020 3613.980 89.260 ;
  LAYER metal3 ;
  RECT 3612.860 86.020 3613.980 89.260 ;
  LAYER metal2 ;
  RECT 3612.860 86.020 3613.980 89.260 ;
  LAYER metal1 ;
  RECT 3612.860 86.020 3613.980 89.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 46.820 3613.980 50.060 ;
  LAYER metal4 ;
  RECT 3612.860 46.820 3613.980 50.060 ;
  LAYER metal3 ;
  RECT 3612.860 46.820 3613.980 50.060 ;
  LAYER metal2 ;
  RECT 3612.860 46.820 3613.980 50.060 ;
  LAYER metal1 ;
  RECT 3612.860 46.820 3613.980 50.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 38.980 3613.980 42.220 ;
  LAYER metal4 ;
  RECT 3612.860 38.980 3613.980 42.220 ;
  LAYER metal3 ;
  RECT 3612.860 38.980 3613.980 42.220 ;
  LAYER metal2 ;
  RECT 3612.860 38.980 3613.980 42.220 ;
  LAYER metal1 ;
  RECT 3612.860 38.980 3613.980 42.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 31.140 3613.980 34.380 ;
  LAYER metal4 ;
  RECT 3612.860 31.140 3613.980 34.380 ;
  LAYER metal3 ;
  RECT 3612.860 31.140 3613.980 34.380 ;
  LAYER metal2 ;
  RECT 3612.860 31.140 3613.980 34.380 ;
  LAYER metal1 ;
  RECT 3612.860 31.140 3613.980 34.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 23.300 3613.980 26.540 ;
  LAYER metal4 ;
  RECT 3612.860 23.300 3613.980 26.540 ;
  LAYER metal3 ;
  RECT 3612.860 23.300 3613.980 26.540 ;
  LAYER metal2 ;
  RECT 3612.860 23.300 3613.980 26.540 ;
  LAYER metal1 ;
  RECT 3612.860 23.300 3613.980 26.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 15.460 3613.980 18.700 ;
  LAYER metal4 ;
  RECT 3612.860 15.460 3613.980 18.700 ;
  LAYER metal3 ;
  RECT 3612.860 15.460 3613.980 18.700 ;
  LAYER metal2 ;
  RECT 3612.860 15.460 3613.980 18.700 ;
  LAYER metal1 ;
  RECT 3612.860 15.460 3613.980 18.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3612.860 7.620 3613.980 10.860 ;
  LAYER metal4 ;
  RECT 3612.860 7.620 3613.980 10.860 ;
  LAYER metal3 ;
  RECT 3612.860 7.620 3613.980 10.860 ;
  LAYER metal2 ;
  RECT 3612.860 7.620 3613.980 10.860 ;
  LAYER metal1 ;
  RECT 3612.860 7.620 3613.980 10.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1693.220 1.120 1696.460 ;
  LAYER metal4 ;
  RECT 0.000 1693.220 1.120 1696.460 ;
  LAYER metal3 ;
  RECT 0.000 1693.220 1.120 1696.460 ;
  LAYER metal2 ;
  RECT 0.000 1693.220 1.120 1696.460 ;
  LAYER metal1 ;
  RECT 0.000 1693.220 1.120 1696.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1685.380 1.120 1688.620 ;
  LAYER metal4 ;
  RECT 0.000 1685.380 1.120 1688.620 ;
  LAYER metal3 ;
  RECT 0.000 1685.380 1.120 1688.620 ;
  LAYER metal2 ;
  RECT 0.000 1685.380 1.120 1688.620 ;
  LAYER metal1 ;
  RECT 0.000 1685.380 1.120 1688.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1677.540 1.120 1680.780 ;
  LAYER metal4 ;
  RECT 0.000 1677.540 1.120 1680.780 ;
  LAYER metal3 ;
  RECT 0.000 1677.540 1.120 1680.780 ;
  LAYER metal2 ;
  RECT 0.000 1677.540 1.120 1680.780 ;
  LAYER metal1 ;
  RECT 0.000 1677.540 1.120 1680.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1669.700 1.120 1672.940 ;
  LAYER metal4 ;
  RECT 0.000 1669.700 1.120 1672.940 ;
  LAYER metal3 ;
  RECT 0.000 1669.700 1.120 1672.940 ;
  LAYER metal2 ;
  RECT 0.000 1669.700 1.120 1672.940 ;
  LAYER metal1 ;
  RECT 0.000 1669.700 1.120 1672.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1661.860 1.120 1665.100 ;
  LAYER metal4 ;
  RECT 0.000 1661.860 1.120 1665.100 ;
  LAYER metal3 ;
  RECT 0.000 1661.860 1.120 1665.100 ;
  LAYER metal2 ;
  RECT 0.000 1661.860 1.120 1665.100 ;
  LAYER metal1 ;
  RECT 0.000 1661.860 1.120 1665.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1654.020 1.120 1657.260 ;
  LAYER metal4 ;
  RECT 0.000 1654.020 1.120 1657.260 ;
  LAYER metal3 ;
  RECT 0.000 1654.020 1.120 1657.260 ;
  LAYER metal2 ;
  RECT 0.000 1654.020 1.120 1657.260 ;
  LAYER metal1 ;
  RECT 0.000 1654.020 1.120 1657.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1614.820 1.120 1618.060 ;
  LAYER metal4 ;
  RECT 0.000 1614.820 1.120 1618.060 ;
  LAYER metal3 ;
  RECT 0.000 1614.820 1.120 1618.060 ;
  LAYER metal2 ;
  RECT 0.000 1614.820 1.120 1618.060 ;
  LAYER metal1 ;
  RECT 0.000 1614.820 1.120 1618.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1606.980 1.120 1610.220 ;
  LAYER metal4 ;
  RECT 0.000 1606.980 1.120 1610.220 ;
  LAYER metal3 ;
  RECT 0.000 1606.980 1.120 1610.220 ;
  LAYER metal2 ;
  RECT 0.000 1606.980 1.120 1610.220 ;
  LAYER metal1 ;
  RECT 0.000 1606.980 1.120 1610.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1599.140 1.120 1602.380 ;
  LAYER metal4 ;
  RECT 0.000 1599.140 1.120 1602.380 ;
  LAYER metal3 ;
  RECT 0.000 1599.140 1.120 1602.380 ;
  LAYER metal2 ;
  RECT 0.000 1599.140 1.120 1602.380 ;
  LAYER metal1 ;
  RECT 0.000 1599.140 1.120 1602.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1591.300 1.120 1594.540 ;
  LAYER metal4 ;
  RECT 0.000 1591.300 1.120 1594.540 ;
  LAYER metal3 ;
  RECT 0.000 1591.300 1.120 1594.540 ;
  LAYER metal2 ;
  RECT 0.000 1591.300 1.120 1594.540 ;
  LAYER metal1 ;
  RECT 0.000 1591.300 1.120 1594.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1583.460 1.120 1586.700 ;
  LAYER metal4 ;
  RECT 0.000 1583.460 1.120 1586.700 ;
  LAYER metal3 ;
  RECT 0.000 1583.460 1.120 1586.700 ;
  LAYER metal2 ;
  RECT 0.000 1583.460 1.120 1586.700 ;
  LAYER metal1 ;
  RECT 0.000 1583.460 1.120 1586.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1575.620 1.120 1578.860 ;
  LAYER metal4 ;
  RECT 0.000 1575.620 1.120 1578.860 ;
  LAYER metal3 ;
  RECT 0.000 1575.620 1.120 1578.860 ;
  LAYER metal2 ;
  RECT 0.000 1575.620 1.120 1578.860 ;
  LAYER metal1 ;
  RECT 0.000 1575.620 1.120 1578.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1536.420 1.120 1539.660 ;
  LAYER metal4 ;
  RECT 0.000 1536.420 1.120 1539.660 ;
  LAYER metal3 ;
  RECT 0.000 1536.420 1.120 1539.660 ;
  LAYER metal2 ;
  RECT 0.000 1536.420 1.120 1539.660 ;
  LAYER metal1 ;
  RECT 0.000 1536.420 1.120 1539.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1528.580 1.120 1531.820 ;
  LAYER metal4 ;
  RECT 0.000 1528.580 1.120 1531.820 ;
  LAYER metal3 ;
  RECT 0.000 1528.580 1.120 1531.820 ;
  LAYER metal2 ;
  RECT 0.000 1528.580 1.120 1531.820 ;
  LAYER metal1 ;
  RECT 0.000 1528.580 1.120 1531.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1520.740 1.120 1523.980 ;
  LAYER metal4 ;
  RECT 0.000 1520.740 1.120 1523.980 ;
  LAYER metal3 ;
  RECT 0.000 1520.740 1.120 1523.980 ;
  LAYER metal2 ;
  RECT 0.000 1520.740 1.120 1523.980 ;
  LAYER metal1 ;
  RECT 0.000 1520.740 1.120 1523.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1512.900 1.120 1516.140 ;
  LAYER metal4 ;
  RECT 0.000 1512.900 1.120 1516.140 ;
  LAYER metal3 ;
  RECT 0.000 1512.900 1.120 1516.140 ;
  LAYER metal2 ;
  RECT 0.000 1512.900 1.120 1516.140 ;
  LAYER metal1 ;
  RECT 0.000 1512.900 1.120 1516.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1505.060 1.120 1508.300 ;
  LAYER metal4 ;
  RECT 0.000 1505.060 1.120 1508.300 ;
  LAYER metal3 ;
  RECT 0.000 1505.060 1.120 1508.300 ;
  LAYER metal2 ;
  RECT 0.000 1505.060 1.120 1508.300 ;
  LAYER metal1 ;
  RECT 0.000 1505.060 1.120 1508.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1497.220 1.120 1500.460 ;
  LAYER metal4 ;
  RECT 0.000 1497.220 1.120 1500.460 ;
  LAYER metal3 ;
  RECT 0.000 1497.220 1.120 1500.460 ;
  LAYER metal2 ;
  RECT 0.000 1497.220 1.120 1500.460 ;
  LAYER metal1 ;
  RECT 0.000 1497.220 1.120 1500.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1458.020 1.120 1461.260 ;
  LAYER metal4 ;
  RECT 0.000 1458.020 1.120 1461.260 ;
  LAYER metal3 ;
  RECT 0.000 1458.020 1.120 1461.260 ;
  LAYER metal2 ;
  RECT 0.000 1458.020 1.120 1461.260 ;
  LAYER metal1 ;
  RECT 0.000 1458.020 1.120 1461.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1450.180 1.120 1453.420 ;
  LAYER metal4 ;
  RECT 0.000 1450.180 1.120 1453.420 ;
  LAYER metal3 ;
  RECT 0.000 1450.180 1.120 1453.420 ;
  LAYER metal2 ;
  RECT 0.000 1450.180 1.120 1453.420 ;
  LAYER metal1 ;
  RECT 0.000 1450.180 1.120 1453.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1442.340 1.120 1445.580 ;
  LAYER metal4 ;
  RECT 0.000 1442.340 1.120 1445.580 ;
  LAYER metal3 ;
  RECT 0.000 1442.340 1.120 1445.580 ;
  LAYER metal2 ;
  RECT 0.000 1442.340 1.120 1445.580 ;
  LAYER metal1 ;
  RECT 0.000 1442.340 1.120 1445.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1434.500 1.120 1437.740 ;
  LAYER metal4 ;
  RECT 0.000 1434.500 1.120 1437.740 ;
  LAYER metal3 ;
  RECT 0.000 1434.500 1.120 1437.740 ;
  LAYER metal2 ;
  RECT 0.000 1434.500 1.120 1437.740 ;
  LAYER metal1 ;
  RECT 0.000 1434.500 1.120 1437.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1426.660 1.120 1429.900 ;
  LAYER metal4 ;
  RECT 0.000 1426.660 1.120 1429.900 ;
  LAYER metal3 ;
  RECT 0.000 1426.660 1.120 1429.900 ;
  LAYER metal2 ;
  RECT 0.000 1426.660 1.120 1429.900 ;
  LAYER metal1 ;
  RECT 0.000 1426.660 1.120 1429.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1418.820 1.120 1422.060 ;
  LAYER metal4 ;
  RECT 0.000 1418.820 1.120 1422.060 ;
  LAYER metal3 ;
  RECT 0.000 1418.820 1.120 1422.060 ;
  LAYER metal2 ;
  RECT 0.000 1418.820 1.120 1422.060 ;
  LAYER metal1 ;
  RECT 0.000 1418.820 1.120 1422.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1379.620 1.120 1382.860 ;
  LAYER metal4 ;
  RECT 0.000 1379.620 1.120 1382.860 ;
  LAYER metal3 ;
  RECT 0.000 1379.620 1.120 1382.860 ;
  LAYER metal2 ;
  RECT 0.000 1379.620 1.120 1382.860 ;
  LAYER metal1 ;
  RECT 0.000 1379.620 1.120 1382.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1371.780 1.120 1375.020 ;
  LAYER metal4 ;
  RECT 0.000 1371.780 1.120 1375.020 ;
  LAYER metal3 ;
  RECT 0.000 1371.780 1.120 1375.020 ;
  LAYER metal2 ;
  RECT 0.000 1371.780 1.120 1375.020 ;
  LAYER metal1 ;
  RECT 0.000 1371.780 1.120 1375.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1363.940 1.120 1367.180 ;
  LAYER metal4 ;
  RECT 0.000 1363.940 1.120 1367.180 ;
  LAYER metal3 ;
  RECT 0.000 1363.940 1.120 1367.180 ;
  LAYER metal2 ;
  RECT 0.000 1363.940 1.120 1367.180 ;
  LAYER metal1 ;
  RECT 0.000 1363.940 1.120 1367.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1356.100 1.120 1359.340 ;
  LAYER metal4 ;
  RECT 0.000 1356.100 1.120 1359.340 ;
  LAYER metal3 ;
  RECT 0.000 1356.100 1.120 1359.340 ;
  LAYER metal2 ;
  RECT 0.000 1356.100 1.120 1359.340 ;
  LAYER metal1 ;
  RECT 0.000 1356.100 1.120 1359.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1348.260 1.120 1351.500 ;
  LAYER metal4 ;
  RECT 0.000 1348.260 1.120 1351.500 ;
  LAYER metal3 ;
  RECT 0.000 1348.260 1.120 1351.500 ;
  LAYER metal2 ;
  RECT 0.000 1348.260 1.120 1351.500 ;
  LAYER metal1 ;
  RECT 0.000 1348.260 1.120 1351.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1340.420 1.120 1343.660 ;
  LAYER metal4 ;
  RECT 0.000 1340.420 1.120 1343.660 ;
  LAYER metal3 ;
  RECT 0.000 1340.420 1.120 1343.660 ;
  LAYER metal2 ;
  RECT 0.000 1340.420 1.120 1343.660 ;
  LAYER metal1 ;
  RECT 0.000 1340.420 1.120 1343.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1301.220 1.120 1304.460 ;
  LAYER metal4 ;
  RECT 0.000 1301.220 1.120 1304.460 ;
  LAYER metal3 ;
  RECT 0.000 1301.220 1.120 1304.460 ;
  LAYER metal2 ;
  RECT 0.000 1301.220 1.120 1304.460 ;
  LAYER metal1 ;
  RECT 0.000 1301.220 1.120 1304.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1293.380 1.120 1296.620 ;
  LAYER metal4 ;
  RECT 0.000 1293.380 1.120 1296.620 ;
  LAYER metal3 ;
  RECT 0.000 1293.380 1.120 1296.620 ;
  LAYER metal2 ;
  RECT 0.000 1293.380 1.120 1296.620 ;
  LAYER metal1 ;
  RECT 0.000 1293.380 1.120 1296.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1285.540 1.120 1288.780 ;
  LAYER metal4 ;
  RECT 0.000 1285.540 1.120 1288.780 ;
  LAYER metal3 ;
  RECT 0.000 1285.540 1.120 1288.780 ;
  LAYER metal2 ;
  RECT 0.000 1285.540 1.120 1288.780 ;
  LAYER metal1 ;
  RECT 0.000 1285.540 1.120 1288.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1277.700 1.120 1280.940 ;
  LAYER metal4 ;
  RECT 0.000 1277.700 1.120 1280.940 ;
  LAYER metal3 ;
  RECT 0.000 1277.700 1.120 1280.940 ;
  LAYER metal2 ;
  RECT 0.000 1277.700 1.120 1280.940 ;
  LAYER metal1 ;
  RECT 0.000 1277.700 1.120 1280.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1269.860 1.120 1273.100 ;
  LAYER metal4 ;
  RECT 0.000 1269.860 1.120 1273.100 ;
  LAYER metal3 ;
  RECT 0.000 1269.860 1.120 1273.100 ;
  LAYER metal2 ;
  RECT 0.000 1269.860 1.120 1273.100 ;
  LAYER metal1 ;
  RECT 0.000 1269.860 1.120 1273.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1262.020 1.120 1265.260 ;
  LAYER metal4 ;
  RECT 0.000 1262.020 1.120 1265.260 ;
  LAYER metal3 ;
  RECT 0.000 1262.020 1.120 1265.260 ;
  LAYER metal2 ;
  RECT 0.000 1262.020 1.120 1265.260 ;
  LAYER metal1 ;
  RECT 0.000 1262.020 1.120 1265.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1222.820 1.120 1226.060 ;
  LAYER metal4 ;
  RECT 0.000 1222.820 1.120 1226.060 ;
  LAYER metal3 ;
  RECT 0.000 1222.820 1.120 1226.060 ;
  LAYER metal2 ;
  RECT 0.000 1222.820 1.120 1226.060 ;
  LAYER metal1 ;
  RECT 0.000 1222.820 1.120 1226.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1214.980 1.120 1218.220 ;
  LAYER metal4 ;
  RECT 0.000 1214.980 1.120 1218.220 ;
  LAYER metal3 ;
  RECT 0.000 1214.980 1.120 1218.220 ;
  LAYER metal2 ;
  RECT 0.000 1214.980 1.120 1218.220 ;
  LAYER metal1 ;
  RECT 0.000 1214.980 1.120 1218.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1207.140 1.120 1210.380 ;
  LAYER metal4 ;
  RECT 0.000 1207.140 1.120 1210.380 ;
  LAYER metal3 ;
  RECT 0.000 1207.140 1.120 1210.380 ;
  LAYER metal2 ;
  RECT 0.000 1207.140 1.120 1210.380 ;
  LAYER metal1 ;
  RECT 0.000 1207.140 1.120 1210.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1199.300 1.120 1202.540 ;
  LAYER metal4 ;
  RECT 0.000 1199.300 1.120 1202.540 ;
  LAYER metal3 ;
  RECT 0.000 1199.300 1.120 1202.540 ;
  LAYER metal2 ;
  RECT 0.000 1199.300 1.120 1202.540 ;
  LAYER metal1 ;
  RECT 0.000 1199.300 1.120 1202.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1191.460 1.120 1194.700 ;
  LAYER metal4 ;
  RECT 0.000 1191.460 1.120 1194.700 ;
  LAYER metal3 ;
  RECT 0.000 1191.460 1.120 1194.700 ;
  LAYER metal2 ;
  RECT 0.000 1191.460 1.120 1194.700 ;
  LAYER metal1 ;
  RECT 0.000 1191.460 1.120 1194.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1183.620 1.120 1186.860 ;
  LAYER metal4 ;
  RECT 0.000 1183.620 1.120 1186.860 ;
  LAYER metal3 ;
  RECT 0.000 1183.620 1.120 1186.860 ;
  LAYER metal2 ;
  RECT 0.000 1183.620 1.120 1186.860 ;
  LAYER metal1 ;
  RECT 0.000 1183.620 1.120 1186.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1144.420 1.120 1147.660 ;
  LAYER metal4 ;
  RECT 0.000 1144.420 1.120 1147.660 ;
  LAYER metal3 ;
  RECT 0.000 1144.420 1.120 1147.660 ;
  LAYER metal2 ;
  RECT 0.000 1144.420 1.120 1147.660 ;
  LAYER metal1 ;
  RECT 0.000 1144.420 1.120 1147.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1136.580 1.120 1139.820 ;
  LAYER metal4 ;
  RECT 0.000 1136.580 1.120 1139.820 ;
  LAYER metal3 ;
  RECT 0.000 1136.580 1.120 1139.820 ;
  LAYER metal2 ;
  RECT 0.000 1136.580 1.120 1139.820 ;
  LAYER metal1 ;
  RECT 0.000 1136.580 1.120 1139.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1128.740 1.120 1131.980 ;
  LAYER metal4 ;
  RECT 0.000 1128.740 1.120 1131.980 ;
  LAYER metal3 ;
  RECT 0.000 1128.740 1.120 1131.980 ;
  LAYER metal2 ;
  RECT 0.000 1128.740 1.120 1131.980 ;
  LAYER metal1 ;
  RECT 0.000 1128.740 1.120 1131.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1120.900 1.120 1124.140 ;
  LAYER metal4 ;
  RECT 0.000 1120.900 1.120 1124.140 ;
  LAYER metal3 ;
  RECT 0.000 1120.900 1.120 1124.140 ;
  LAYER metal2 ;
  RECT 0.000 1120.900 1.120 1124.140 ;
  LAYER metal1 ;
  RECT 0.000 1120.900 1.120 1124.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1113.060 1.120 1116.300 ;
  LAYER metal4 ;
  RECT 0.000 1113.060 1.120 1116.300 ;
  LAYER metal3 ;
  RECT 0.000 1113.060 1.120 1116.300 ;
  LAYER metal2 ;
  RECT 0.000 1113.060 1.120 1116.300 ;
  LAYER metal1 ;
  RECT 0.000 1113.060 1.120 1116.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1105.220 1.120 1108.460 ;
  LAYER metal4 ;
  RECT 0.000 1105.220 1.120 1108.460 ;
  LAYER metal3 ;
  RECT 0.000 1105.220 1.120 1108.460 ;
  LAYER metal2 ;
  RECT 0.000 1105.220 1.120 1108.460 ;
  LAYER metal1 ;
  RECT 0.000 1105.220 1.120 1108.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1066.020 1.120 1069.260 ;
  LAYER metal4 ;
  RECT 0.000 1066.020 1.120 1069.260 ;
  LAYER metal3 ;
  RECT 0.000 1066.020 1.120 1069.260 ;
  LAYER metal2 ;
  RECT 0.000 1066.020 1.120 1069.260 ;
  LAYER metal1 ;
  RECT 0.000 1066.020 1.120 1069.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1058.180 1.120 1061.420 ;
  LAYER metal4 ;
  RECT 0.000 1058.180 1.120 1061.420 ;
  LAYER metal3 ;
  RECT 0.000 1058.180 1.120 1061.420 ;
  LAYER metal2 ;
  RECT 0.000 1058.180 1.120 1061.420 ;
  LAYER metal1 ;
  RECT 0.000 1058.180 1.120 1061.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1050.340 1.120 1053.580 ;
  LAYER metal4 ;
  RECT 0.000 1050.340 1.120 1053.580 ;
  LAYER metal3 ;
  RECT 0.000 1050.340 1.120 1053.580 ;
  LAYER metal2 ;
  RECT 0.000 1050.340 1.120 1053.580 ;
  LAYER metal1 ;
  RECT 0.000 1050.340 1.120 1053.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1042.500 1.120 1045.740 ;
  LAYER metal4 ;
  RECT 0.000 1042.500 1.120 1045.740 ;
  LAYER metal3 ;
  RECT 0.000 1042.500 1.120 1045.740 ;
  LAYER metal2 ;
  RECT 0.000 1042.500 1.120 1045.740 ;
  LAYER metal1 ;
  RECT 0.000 1042.500 1.120 1045.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1034.660 1.120 1037.900 ;
  LAYER metal4 ;
  RECT 0.000 1034.660 1.120 1037.900 ;
  LAYER metal3 ;
  RECT 0.000 1034.660 1.120 1037.900 ;
  LAYER metal2 ;
  RECT 0.000 1034.660 1.120 1037.900 ;
  LAYER metal1 ;
  RECT 0.000 1034.660 1.120 1037.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 1026.820 1.120 1030.060 ;
  LAYER metal4 ;
  RECT 0.000 1026.820 1.120 1030.060 ;
  LAYER metal3 ;
  RECT 0.000 1026.820 1.120 1030.060 ;
  LAYER metal2 ;
  RECT 0.000 1026.820 1.120 1030.060 ;
  LAYER metal1 ;
  RECT 0.000 1026.820 1.120 1030.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 987.620 1.120 990.860 ;
  LAYER metal4 ;
  RECT 0.000 987.620 1.120 990.860 ;
  LAYER metal3 ;
  RECT 0.000 987.620 1.120 990.860 ;
  LAYER metal2 ;
  RECT 0.000 987.620 1.120 990.860 ;
  LAYER metal1 ;
  RECT 0.000 987.620 1.120 990.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 979.780 1.120 983.020 ;
  LAYER metal4 ;
  RECT 0.000 979.780 1.120 983.020 ;
  LAYER metal3 ;
  RECT 0.000 979.780 1.120 983.020 ;
  LAYER metal2 ;
  RECT 0.000 979.780 1.120 983.020 ;
  LAYER metal1 ;
  RECT 0.000 979.780 1.120 983.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 971.940 1.120 975.180 ;
  LAYER metal4 ;
  RECT 0.000 971.940 1.120 975.180 ;
  LAYER metal3 ;
  RECT 0.000 971.940 1.120 975.180 ;
  LAYER metal2 ;
  RECT 0.000 971.940 1.120 975.180 ;
  LAYER metal1 ;
  RECT 0.000 971.940 1.120 975.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 964.100 1.120 967.340 ;
  LAYER metal4 ;
  RECT 0.000 964.100 1.120 967.340 ;
  LAYER metal3 ;
  RECT 0.000 964.100 1.120 967.340 ;
  LAYER metal2 ;
  RECT 0.000 964.100 1.120 967.340 ;
  LAYER metal1 ;
  RECT 0.000 964.100 1.120 967.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 956.260 1.120 959.500 ;
  LAYER metal4 ;
  RECT 0.000 956.260 1.120 959.500 ;
  LAYER metal3 ;
  RECT 0.000 956.260 1.120 959.500 ;
  LAYER metal2 ;
  RECT 0.000 956.260 1.120 959.500 ;
  LAYER metal1 ;
  RECT 0.000 956.260 1.120 959.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 948.420 1.120 951.660 ;
  LAYER metal4 ;
  RECT 0.000 948.420 1.120 951.660 ;
  LAYER metal3 ;
  RECT 0.000 948.420 1.120 951.660 ;
  LAYER metal2 ;
  RECT 0.000 948.420 1.120 951.660 ;
  LAYER metal1 ;
  RECT 0.000 948.420 1.120 951.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 909.220 1.120 912.460 ;
  LAYER metal4 ;
  RECT 0.000 909.220 1.120 912.460 ;
  LAYER metal3 ;
  RECT 0.000 909.220 1.120 912.460 ;
  LAYER metal2 ;
  RECT 0.000 909.220 1.120 912.460 ;
  LAYER metal1 ;
  RECT 0.000 909.220 1.120 912.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 901.380 1.120 904.620 ;
  LAYER metal4 ;
  RECT 0.000 901.380 1.120 904.620 ;
  LAYER metal3 ;
  RECT 0.000 901.380 1.120 904.620 ;
  LAYER metal2 ;
  RECT 0.000 901.380 1.120 904.620 ;
  LAYER metal1 ;
  RECT 0.000 901.380 1.120 904.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 893.540 1.120 896.780 ;
  LAYER metal4 ;
  RECT 0.000 893.540 1.120 896.780 ;
  LAYER metal3 ;
  RECT 0.000 893.540 1.120 896.780 ;
  LAYER metal2 ;
  RECT 0.000 893.540 1.120 896.780 ;
  LAYER metal1 ;
  RECT 0.000 893.540 1.120 896.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 885.700 1.120 888.940 ;
  LAYER metal4 ;
  RECT 0.000 885.700 1.120 888.940 ;
  LAYER metal3 ;
  RECT 0.000 885.700 1.120 888.940 ;
  LAYER metal2 ;
  RECT 0.000 885.700 1.120 888.940 ;
  LAYER metal1 ;
  RECT 0.000 885.700 1.120 888.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 877.860 1.120 881.100 ;
  LAYER metal4 ;
  RECT 0.000 877.860 1.120 881.100 ;
  LAYER metal3 ;
  RECT 0.000 877.860 1.120 881.100 ;
  LAYER metal2 ;
  RECT 0.000 877.860 1.120 881.100 ;
  LAYER metal1 ;
  RECT 0.000 877.860 1.120 881.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 870.020 1.120 873.260 ;
  LAYER metal4 ;
  RECT 0.000 870.020 1.120 873.260 ;
  LAYER metal3 ;
  RECT 0.000 870.020 1.120 873.260 ;
  LAYER metal2 ;
  RECT 0.000 870.020 1.120 873.260 ;
  LAYER metal1 ;
  RECT 0.000 870.020 1.120 873.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 830.820 1.120 834.060 ;
  LAYER metal4 ;
  RECT 0.000 830.820 1.120 834.060 ;
  LAYER metal3 ;
  RECT 0.000 830.820 1.120 834.060 ;
  LAYER metal2 ;
  RECT 0.000 830.820 1.120 834.060 ;
  LAYER metal1 ;
  RECT 0.000 830.820 1.120 834.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 822.980 1.120 826.220 ;
  LAYER metal4 ;
  RECT 0.000 822.980 1.120 826.220 ;
  LAYER metal3 ;
  RECT 0.000 822.980 1.120 826.220 ;
  LAYER metal2 ;
  RECT 0.000 822.980 1.120 826.220 ;
  LAYER metal1 ;
  RECT 0.000 822.980 1.120 826.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 815.140 1.120 818.380 ;
  LAYER metal4 ;
  RECT 0.000 815.140 1.120 818.380 ;
  LAYER metal3 ;
  RECT 0.000 815.140 1.120 818.380 ;
  LAYER metal2 ;
  RECT 0.000 815.140 1.120 818.380 ;
  LAYER metal1 ;
  RECT 0.000 815.140 1.120 818.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 807.300 1.120 810.540 ;
  LAYER metal4 ;
  RECT 0.000 807.300 1.120 810.540 ;
  LAYER metal3 ;
  RECT 0.000 807.300 1.120 810.540 ;
  LAYER metal2 ;
  RECT 0.000 807.300 1.120 810.540 ;
  LAYER metal1 ;
  RECT 0.000 807.300 1.120 810.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 799.460 1.120 802.700 ;
  LAYER metal4 ;
  RECT 0.000 799.460 1.120 802.700 ;
  LAYER metal3 ;
  RECT 0.000 799.460 1.120 802.700 ;
  LAYER metal2 ;
  RECT 0.000 799.460 1.120 802.700 ;
  LAYER metal1 ;
  RECT 0.000 799.460 1.120 802.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 791.620 1.120 794.860 ;
  LAYER metal4 ;
  RECT 0.000 791.620 1.120 794.860 ;
  LAYER metal3 ;
  RECT 0.000 791.620 1.120 794.860 ;
  LAYER metal2 ;
  RECT 0.000 791.620 1.120 794.860 ;
  LAYER metal1 ;
  RECT 0.000 791.620 1.120 794.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 752.420 1.120 755.660 ;
  LAYER metal4 ;
  RECT 0.000 752.420 1.120 755.660 ;
  LAYER metal3 ;
  RECT 0.000 752.420 1.120 755.660 ;
  LAYER metal2 ;
  RECT 0.000 752.420 1.120 755.660 ;
  LAYER metal1 ;
  RECT 0.000 752.420 1.120 755.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 744.580 1.120 747.820 ;
  LAYER metal4 ;
  RECT 0.000 744.580 1.120 747.820 ;
  LAYER metal3 ;
  RECT 0.000 744.580 1.120 747.820 ;
  LAYER metal2 ;
  RECT 0.000 744.580 1.120 747.820 ;
  LAYER metal1 ;
  RECT 0.000 744.580 1.120 747.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 736.740 1.120 739.980 ;
  LAYER metal4 ;
  RECT 0.000 736.740 1.120 739.980 ;
  LAYER metal3 ;
  RECT 0.000 736.740 1.120 739.980 ;
  LAYER metal2 ;
  RECT 0.000 736.740 1.120 739.980 ;
  LAYER metal1 ;
  RECT 0.000 736.740 1.120 739.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 728.900 1.120 732.140 ;
  LAYER metal4 ;
  RECT 0.000 728.900 1.120 732.140 ;
  LAYER metal3 ;
  RECT 0.000 728.900 1.120 732.140 ;
  LAYER metal2 ;
  RECT 0.000 728.900 1.120 732.140 ;
  LAYER metal1 ;
  RECT 0.000 728.900 1.120 732.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 721.060 1.120 724.300 ;
  LAYER metal4 ;
  RECT 0.000 721.060 1.120 724.300 ;
  LAYER metal3 ;
  RECT 0.000 721.060 1.120 724.300 ;
  LAYER metal2 ;
  RECT 0.000 721.060 1.120 724.300 ;
  LAYER metal1 ;
  RECT 0.000 721.060 1.120 724.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 713.220 1.120 716.460 ;
  LAYER metal4 ;
  RECT 0.000 713.220 1.120 716.460 ;
  LAYER metal3 ;
  RECT 0.000 713.220 1.120 716.460 ;
  LAYER metal2 ;
  RECT 0.000 713.220 1.120 716.460 ;
  LAYER metal1 ;
  RECT 0.000 713.220 1.120 716.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 674.020 1.120 677.260 ;
  LAYER metal4 ;
  RECT 0.000 674.020 1.120 677.260 ;
  LAYER metal3 ;
  RECT 0.000 674.020 1.120 677.260 ;
  LAYER metal2 ;
  RECT 0.000 674.020 1.120 677.260 ;
  LAYER metal1 ;
  RECT 0.000 674.020 1.120 677.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 666.180 1.120 669.420 ;
  LAYER metal4 ;
  RECT 0.000 666.180 1.120 669.420 ;
  LAYER metal3 ;
  RECT 0.000 666.180 1.120 669.420 ;
  LAYER metal2 ;
  RECT 0.000 666.180 1.120 669.420 ;
  LAYER metal1 ;
  RECT 0.000 666.180 1.120 669.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 658.340 1.120 661.580 ;
  LAYER metal4 ;
  RECT 0.000 658.340 1.120 661.580 ;
  LAYER metal3 ;
  RECT 0.000 658.340 1.120 661.580 ;
  LAYER metal2 ;
  RECT 0.000 658.340 1.120 661.580 ;
  LAYER metal1 ;
  RECT 0.000 658.340 1.120 661.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 650.500 1.120 653.740 ;
  LAYER metal4 ;
  RECT 0.000 650.500 1.120 653.740 ;
  LAYER metal3 ;
  RECT 0.000 650.500 1.120 653.740 ;
  LAYER metal2 ;
  RECT 0.000 650.500 1.120 653.740 ;
  LAYER metal1 ;
  RECT 0.000 650.500 1.120 653.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 642.660 1.120 645.900 ;
  LAYER metal4 ;
  RECT 0.000 642.660 1.120 645.900 ;
  LAYER metal3 ;
  RECT 0.000 642.660 1.120 645.900 ;
  LAYER metal2 ;
  RECT 0.000 642.660 1.120 645.900 ;
  LAYER metal1 ;
  RECT 0.000 642.660 1.120 645.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 634.820 1.120 638.060 ;
  LAYER metal4 ;
  RECT 0.000 634.820 1.120 638.060 ;
  LAYER metal3 ;
  RECT 0.000 634.820 1.120 638.060 ;
  LAYER metal2 ;
  RECT 0.000 634.820 1.120 638.060 ;
  LAYER metal1 ;
  RECT 0.000 634.820 1.120 638.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 595.620 1.120 598.860 ;
  LAYER metal4 ;
  RECT 0.000 595.620 1.120 598.860 ;
  LAYER metal3 ;
  RECT 0.000 595.620 1.120 598.860 ;
  LAYER metal2 ;
  RECT 0.000 595.620 1.120 598.860 ;
  LAYER metal1 ;
  RECT 0.000 595.620 1.120 598.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 587.780 1.120 591.020 ;
  LAYER metal4 ;
  RECT 0.000 587.780 1.120 591.020 ;
  LAYER metal3 ;
  RECT 0.000 587.780 1.120 591.020 ;
  LAYER metal2 ;
  RECT 0.000 587.780 1.120 591.020 ;
  LAYER metal1 ;
  RECT 0.000 587.780 1.120 591.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 579.940 1.120 583.180 ;
  LAYER metal4 ;
  RECT 0.000 579.940 1.120 583.180 ;
  LAYER metal3 ;
  RECT 0.000 579.940 1.120 583.180 ;
  LAYER metal2 ;
  RECT 0.000 579.940 1.120 583.180 ;
  LAYER metal1 ;
  RECT 0.000 579.940 1.120 583.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 572.100 1.120 575.340 ;
  LAYER metal4 ;
  RECT 0.000 572.100 1.120 575.340 ;
  LAYER metal3 ;
  RECT 0.000 572.100 1.120 575.340 ;
  LAYER metal2 ;
  RECT 0.000 572.100 1.120 575.340 ;
  LAYER metal1 ;
  RECT 0.000 572.100 1.120 575.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 564.260 1.120 567.500 ;
  LAYER metal4 ;
  RECT 0.000 564.260 1.120 567.500 ;
  LAYER metal3 ;
  RECT 0.000 564.260 1.120 567.500 ;
  LAYER metal2 ;
  RECT 0.000 564.260 1.120 567.500 ;
  LAYER metal1 ;
  RECT 0.000 564.260 1.120 567.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 556.420 1.120 559.660 ;
  LAYER metal4 ;
  RECT 0.000 556.420 1.120 559.660 ;
  LAYER metal3 ;
  RECT 0.000 556.420 1.120 559.660 ;
  LAYER metal2 ;
  RECT 0.000 556.420 1.120 559.660 ;
  LAYER metal1 ;
  RECT 0.000 556.420 1.120 559.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 517.220 1.120 520.460 ;
  LAYER metal4 ;
  RECT 0.000 517.220 1.120 520.460 ;
  LAYER metal3 ;
  RECT 0.000 517.220 1.120 520.460 ;
  LAYER metal2 ;
  RECT 0.000 517.220 1.120 520.460 ;
  LAYER metal1 ;
  RECT 0.000 517.220 1.120 520.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 509.380 1.120 512.620 ;
  LAYER metal4 ;
  RECT 0.000 509.380 1.120 512.620 ;
  LAYER metal3 ;
  RECT 0.000 509.380 1.120 512.620 ;
  LAYER metal2 ;
  RECT 0.000 509.380 1.120 512.620 ;
  LAYER metal1 ;
  RECT 0.000 509.380 1.120 512.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 501.540 1.120 504.780 ;
  LAYER metal4 ;
  RECT 0.000 501.540 1.120 504.780 ;
  LAYER metal3 ;
  RECT 0.000 501.540 1.120 504.780 ;
  LAYER metal2 ;
  RECT 0.000 501.540 1.120 504.780 ;
  LAYER metal1 ;
  RECT 0.000 501.540 1.120 504.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 493.700 1.120 496.940 ;
  LAYER metal4 ;
  RECT 0.000 493.700 1.120 496.940 ;
  LAYER metal3 ;
  RECT 0.000 493.700 1.120 496.940 ;
  LAYER metal2 ;
  RECT 0.000 493.700 1.120 496.940 ;
  LAYER metal1 ;
  RECT 0.000 493.700 1.120 496.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 485.860 1.120 489.100 ;
  LAYER metal4 ;
  RECT 0.000 485.860 1.120 489.100 ;
  LAYER metal3 ;
  RECT 0.000 485.860 1.120 489.100 ;
  LAYER metal2 ;
  RECT 0.000 485.860 1.120 489.100 ;
  LAYER metal1 ;
  RECT 0.000 485.860 1.120 489.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 478.020 1.120 481.260 ;
  LAYER metal4 ;
  RECT 0.000 478.020 1.120 481.260 ;
  LAYER metal3 ;
  RECT 0.000 478.020 1.120 481.260 ;
  LAYER metal2 ;
  RECT 0.000 478.020 1.120 481.260 ;
  LAYER metal1 ;
  RECT 0.000 478.020 1.120 481.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 438.820 1.120 442.060 ;
  LAYER metal4 ;
  RECT 0.000 438.820 1.120 442.060 ;
  LAYER metal3 ;
  RECT 0.000 438.820 1.120 442.060 ;
  LAYER metal2 ;
  RECT 0.000 438.820 1.120 442.060 ;
  LAYER metal1 ;
  RECT 0.000 438.820 1.120 442.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 430.980 1.120 434.220 ;
  LAYER metal4 ;
  RECT 0.000 430.980 1.120 434.220 ;
  LAYER metal3 ;
  RECT 0.000 430.980 1.120 434.220 ;
  LAYER metal2 ;
  RECT 0.000 430.980 1.120 434.220 ;
  LAYER metal1 ;
  RECT 0.000 430.980 1.120 434.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 423.140 1.120 426.380 ;
  LAYER metal4 ;
  RECT 0.000 423.140 1.120 426.380 ;
  LAYER metal3 ;
  RECT 0.000 423.140 1.120 426.380 ;
  LAYER metal2 ;
  RECT 0.000 423.140 1.120 426.380 ;
  LAYER metal1 ;
  RECT 0.000 423.140 1.120 426.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 415.300 1.120 418.540 ;
  LAYER metal4 ;
  RECT 0.000 415.300 1.120 418.540 ;
  LAYER metal3 ;
  RECT 0.000 415.300 1.120 418.540 ;
  LAYER metal2 ;
  RECT 0.000 415.300 1.120 418.540 ;
  LAYER metal1 ;
  RECT 0.000 415.300 1.120 418.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 407.460 1.120 410.700 ;
  LAYER metal4 ;
  RECT 0.000 407.460 1.120 410.700 ;
  LAYER metal3 ;
  RECT 0.000 407.460 1.120 410.700 ;
  LAYER metal2 ;
  RECT 0.000 407.460 1.120 410.700 ;
  LAYER metal1 ;
  RECT 0.000 407.460 1.120 410.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 399.620 1.120 402.860 ;
  LAYER metal4 ;
  RECT 0.000 399.620 1.120 402.860 ;
  LAYER metal3 ;
  RECT 0.000 399.620 1.120 402.860 ;
  LAYER metal2 ;
  RECT 0.000 399.620 1.120 402.860 ;
  LAYER metal1 ;
  RECT 0.000 399.620 1.120 402.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 360.420 1.120 363.660 ;
  LAYER metal4 ;
  RECT 0.000 360.420 1.120 363.660 ;
  LAYER metal3 ;
  RECT 0.000 360.420 1.120 363.660 ;
  LAYER metal2 ;
  RECT 0.000 360.420 1.120 363.660 ;
  LAYER metal1 ;
  RECT 0.000 360.420 1.120 363.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 352.580 1.120 355.820 ;
  LAYER metal4 ;
  RECT 0.000 352.580 1.120 355.820 ;
  LAYER metal3 ;
  RECT 0.000 352.580 1.120 355.820 ;
  LAYER metal2 ;
  RECT 0.000 352.580 1.120 355.820 ;
  LAYER metal1 ;
  RECT 0.000 352.580 1.120 355.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 344.740 1.120 347.980 ;
  LAYER metal4 ;
  RECT 0.000 344.740 1.120 347.980 ;
  LAYER metal3 ;
  RECT 0.000 344.740 1.120 347.980 ;
  LAYER metal2 ;
  RECT 0.000 344.740 1.120 347.980 ;
  LAYER metal1 ;
  RECT 0.000 344.740 1.120 347.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 336.900 1.120 340.140 ;
  LAYER metal4 ;
  RECT 0.000 336.900 1.120 340.140 ;
  LAYER metal3 ;
  RECT 0.000 336.900 1.120 340.140 ;
  LAYER metal2 ;
  RECT 0.000 336.900 1.120 340.140 ;
  LAYER metal1 ;
  RECT 0.000 336.900 1.120 340.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 329.060 1.120 332.300 ;
  LAYER metal4 ;
  RECT 0.000 329.060 1.120 332.300 ;
  LAYER metal3 ;
  RECT 0.000 329.060 1.120 332.300 ;
  LAYER metal2 ;
  RECT 0.000 329.060 1.120 332.300 ;
  LAYER metal1 ;
  RECT 0.000 329.060 1.120 332.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 321.220 1.120 324.460 ;
  LAYER metal4 ;
  RECT 0.000 321.220 1.120 324.460 ;
  LAYER metal3 ;
  RECT 0.000 321.220 1.120 324.460 ;
  LAYER metal2 ;
  RECT 0.000 321.220 1.120 324.460 ;
  LAYER metal1 ;
  RECT 0.000 321.220 1.120 324.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 282.020 1.120 285.260 ;
  LAYER metal4 ;
  RECT 0.000 282.020 1.120 285.260 ;
  LAYER metal3 ;
  RECT 0.000 282.020 1.120 285.260 ;
  LAYER metal2 ;
  RECT 0.000 282.020 1.120 285.260 ;
  LAYER metal1 ;
  RECT 0.000 282.020 1.120 285.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 274.180 1.120 277.420 ;
  LAYER metal4 ;
  RECT 0.000 274.180 1.120 277.420 ;
  LAYER metal3 ;
  RECT 0.000 274.180 1.120 277.420 ;
  LAYER metal2 ;
  RECT 0.000 274.180 1.120 277.420 ;
  LAYER metal1 ;
  RECT 0.000 274.180 1.120 277.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 266.340 1.120 269.580 ;
  LAYER metal4 ;
  RECT 0.000 266.340 1.120 269.580 ;
  LAYER metal3 ;
  RECT 0.000 266.340 1.120 269.580 ;
  LAYER metal2 ;
  RECT 0.000 266.340 1.120 269.580 ;
  LAYER metal1 ;
  RECT 0.000 266.340 1.120 269.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 258.500 1.120 261.740 ;
  LAYER metal4 ;
  RECT 0.000 258.500 1.120 261.740 ;
  LAYER metal3 ;
  RECT 0.000 258.500 1.120 261.740 ;
  LAYER metal2 ;
  RECT 0.000 258.500 1.120 261.740 ;
  LAYER metal1 ;
  RECT 0.000 258.500 1.120 261.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 250.660 1.120 253.900 ;
  LAYER metal4 ;
  RECT 0.000 250.660 1.120 253.900 ;
  LAYER metal3 ;
  RECT 0.000 250.660 1.120 253.900 ;
  LAYER metal2 ;
  RECT 0.000 250.660 1.120 253.900 ;
  LAYER metal1 ;
  RECT 0.000 250.660 1.120 253.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 242.820 1.120 246.060 ;
  LAYER metal4 ;
  RECT 0.000 242.820 1.120 246.060 ;
  LAYER metal3 ;
  RECT 0.000 242.820 1.120 246.060 ;
  LAYER metal2 ;
  RECT 0.000 242.820 1.120 246.060 ;
  LAYER metal1 ;
  RECT 0.000 242.820 1.120 246.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 203.620 1.120 206.860 ;
  LAYER metal4 ;
  RECT 0.000 203.620 1.120 206.860 ;
  LAYER metal3 ;
  RECT 0.000 203.620 1.120 206.860 ;
  LAYER metal2 ;
  RECT 0.000 203.620 1.120 206.860 ;
  LAYER metal1 ;
  RECT 0.000 203.620 1.120 206.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER metal4 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER metal3 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER metal2 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER metal1 ;
  RECT 0.000 195.780 1.120 199.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER metal4 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER metal3 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER metal2 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER metal1 ;
  RECT 0.000 187.940 1.120 191.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER metal4 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER metal3 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER metal2 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER metal1 ;
  RECT 0.000 180.100 1.120 183.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER metal4 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER metal3 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER metal2 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER metal1 ;
  RECT 0.000 172.260 1.120 175.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER metal4 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER metal3 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER metal2 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER metal1 ;
  RECT 0.000 164.420 1.120 167.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER metal4 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER metal3 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER metal2 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER metal1 ;
  RECT 0.000 125.220 1.120 128.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER metal4 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER metal3 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER metal2 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER metal1 ;
  RECT 0.000 117.380 1.120 120.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER metal4 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER metal3 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER metal2 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER metal1 ;
  RECT 0.000 109.540 1.120 112.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER metal4 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER metal3 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER metal2 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER metal1 ;
  RECT 0.000 101.700 1.120 104.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER metal4 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER metal3 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER metal2 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER metal1 ;
  RECT 0.000 93.860 1.120 97.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER metal4 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER metal3 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER metal2 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER metal1 ;
  RECT 0.000 86.020 1.120 89.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER metal4 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER metal3 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER metal2 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER metal1 ;
  RECT 0.000 46.820 1.120 50.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER metal4 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER metal3 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER metal2 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER metal1 ;
  RECT 0.000 38.980 1.120 42.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER metal4 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER metal3 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER metal2 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER metal1 ;
  RECT 0.000 31.140 1.120 34.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER metal4 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER metal3 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER metal2 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER metal1 ;
  RECT 0.000 23.300 1.120 26.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER metal4 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER metal3 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER metal2 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER metal1 ;
  RECT 0.000 15.460 1.120 18.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER metal4 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER metal3 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER metal2 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER metal1 ;
  RECT 0.000 7.620 1.120 10.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3587.720 1710.800 3591.260 1711.920 ;
  LAYER metal4 ;
  RECT 3587.720 1710.800 3591.260 1711.920 ;
  LAYER metal3 ;
  RECT 3587.720 1710.800 3591.260 1711.920 ;
  LAYER metal2 ;
  RECT 3587.720 1710.800 3591.260 1711.920 ;
  LAYER metal1 ;
  RECT 3587.720 1710.800 3591.260 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3579.040 1710.800 3582.580 1711.920 ;
  LAYER metal4 ;
  RECT 3579.040 1710.800 3582.580 1711.920 ;
  LAYER metal3 ;
  RECT 3579.040 1710.800 3582.580 1711.920 ;
  LAYER metal2 ;
  RECT 3579.040 1710.800 3582.580 1711.920 ;
  LAYER metal1 ;
  RECT 3579.040 1710.800 3582.580 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.360 1710.800 3573.900 1711.920 ;
  LAYER metal4 ;
  RECT 3570.360 1710.800 3573.900 1711.920 ;
  LAYER metal3 ;
  RECT 3570.360 1710.800 3573.900 1711.920 ;
  LAYER metal2 ;
  RECT 3570.360 1710.800 3573.900 1711.920 ;
  LAYER metal1 ;
  RECT 3570.360 1710.800 3573.900 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3561.680 1710.800 3565.220 1711.920 ;
  LAYER metal4 ;
  RECT 3561.680 1710.800 3565.220 1711.920 ;
  LAYER metal3 ;
  RECT 3561.680 1710.800 3565.220 1711.920 ;
  LAYER metal2 ;
  RECT 3561.680 1710.800 3565.220 1711.920 ;
  LAYER metal1 ;
  RECT 3561.680 1710.800 3565.220 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3553.000 1710.800 3556.540 1711.920 ;
  LAYER metal4 ;
  RECT 3553.000 1710.800 3556.540 1711.920 ;
  LAYER metal3 ;
  RECT 3553.000 1710.800 3556.540 1711.920 ;
  LAYER metal2 ;
  RECT 3553.000 1710.800 3556.540 1711.920 ;
  LAYER metal1 ;
  RECT 3553.000 1710.800 3556.540 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3544.320 1710.800 3547.860 1711.920 ;
  LAYER metal4 ;
  RECT 3544.320 1710.800 3547.860 1711.920 ;
  LAYER metal3 ;
  RECT 3544.320 1710.800 3547.860 1711.920 ;
  LAYER metal2 ;
  RECT 3544.320 1710.800 3547.860 1711.920 ;
  LAYER metal1 ;
  RECT 3544.320 1710.800 3547.860 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3500.920 1710.800 3504.460 1711.920 ;
  LAYER metal4 ;
  RECT 3500.920 1710.800 3504.460 1711.920 ;
  LAYER metal3 ;
  RECT 3500.920 1710.800 3504.460 1711.920 ;
  LAYER metal2 ;
  RECT 3500.920 1710.800 3504.460 1711.920 ;
  LAYER metal1 ;
  RECT 3500.920 1710.800 3504.460 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3492.240 1710.800 3495.780 1711.920 ;
  LAYER metal4 ;
  RECT 3492.240 1710.800 3495.780 1711.920 ;
  LAYER metal3 ;
  RECT 3492.240 1710.800 3495.780 1711.920 ;
  LAYER metal2 ;
  RECT 3492.240 1710.800 3495.780 1711.920 ;
  LAYER metal1 ;
  RECT 3492.240 1710.800 3495.780 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3483.560 1710.800 3487.100 1711.920 ;
  LAYER metal4 ;
  RECT 3483.560 1710.800 3487.100 1711.920 ;
  LAYER metal3 ;
  RECT 3483.560 1710.800 3487.100 1711.920 ;
  LAYER metal2 ;
  RECT 3483.560 1710.800 3487.100 1711.920 ;
  LAYER metal1 ;
  RECT 3483.560 1710.800 3487.100 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3474.880 1710.800 3478.420 1711.920 ;
  LAYER metal4 ;
  RECT 3474.880 1710.800 3478.420 1711.920 ;
  LAYER metal3 ;
  RECT 3474.880 1710.800 3478.420 1711.920 ;
  LAYER metal2 ;
  RECT 3474.880 1710.800 3478.420 1711.920 ;
  LAYER metal1 ;
  RECT 3474.880 1710.800 3478.420 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3466.200 1710.800 3469.740 1711.920 ;
  LAYER metal4 ;
  RECT 3466.200 1710.800 3469.740 1711.920 ;
  LAYER metal3 ;
  RECT 3466.200 1710.800 3469.740 1711.920 ;
  LAYER metal2 ;
  RECT 3466.200 1710.800 3469.740 1711.920 ;
  LAYER metal1 ;
  RECT 3466.200 1710.800 3469.740 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3457.520 1710.800 3461.060 1711.920 ;
  LAYER metal4 ;
  RECT 3457.520 1710.800 3461.060 1711.920 ;
  LAYER metal3 ;
  RECT 3457.520 1710.800 3461.060 1711.920 ;
  LAYER metal2 ;
  RECT 3457.520 1710.800 3461.060 1711.920 ;
  LAYER metal1 ;
  RECT 3457.520 1710.800 3461.060 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3414.120 1710.800 3417.660 1711.920 ;
  LAYER metal4 ;
  RECT 3414.120 1710.800 3417.660 1711.920 ;
  LAYER metal3 ;
  RECT 3414.120 1710.800 3417.660 1711.920 ;
  LAYER metal2 ;
  RECT 3414.120 1710.800 3417.660 1711.920 ;
  LAYER metal1 ;
  RECT 3414.120 1710.800 3417.660 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3405.440 1710.800 3408.980 1711.920 ;
  LAYER metal4 ;
  RECT 3405.440 1710.800 3408.980 1711.920 ;
  LAYER metal3 ;
  RECT 3405.440 1710.800 3408.980 1711.920 ;
  LAYER metal2 ;
  RECT 3405.440 1710.800 3408.980 1711.920 ;
  LAYER metal1 ;
  RECT 3405.440 1710.800 3408.980 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3396.760 1710.800 3400.300 1711.920 ;
  LAYER metal4 ;
  RECT 3396.760 1710.800 3400.300 1711.920 ;
  LAYER metal3 ;
  RECT 3396.760 1710.800 3400.300 1711.920 ;
  LAYER metal2 ;
  RECT 3396.760 1710.800 3400.300 1711.920 ;
  LAYER metal1 ;
  RECT 3396.760 1710.800 3400.300 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3388.080 1710.800 3391.620 1711.920 ;
  LAYER metal4 ;
  RECT 3388.080 1710.800 3391.620 1711.920 ;
  LAYER metal3 ;
  RECT 3388.080 1710.800 3391.620 1711.920 ;
  LAYER metal2 ;
  RECT 3388.080 1710.800 3391.620 1711.920 ;
  LAYER metal1 ;
  RECT 3388.080 1710.800 3391.620 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3379.400 1710.800 3382.940 1711.920 ;
  LAYER metal4 ;
  RECT 3379.400 1710.800 3382.940 1711.920 ;
  LAYER metal3 ;
  RECT 3379.400 1710.800 3382.940 1711.920 ;
  LAYER metal2 ;
  RECT 3379.400 1710.800 3382.940 1711.920 ;
  LAYER metal1 ;
  RECT 3379.400 1710.800 3382.940 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3370.720 1710.800 3374.260 1711.920 ;
  LAYER metal4 ;
  RECT 3370.720 1710.800 3374.260 1711.920 ;
  LAYER metal3 ;
  RECT 3370.720 1710.800 3374.260 1711.920 ;
  LAYER metal2 ;
  RECT 3370.720 1710.800 3374.260 1711.920 ;
  LAYER metal1 ;
  RECT 3370.720 1710.800 3374.260 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3327.320 1710.800 3330.860 1711.920 ;
  LAYER metal4 ;
  RECT 3327.320 1710.800 3330.860 1711.920 ;
  LAYER metal3 ;
  RECT 3327.320 1710.800 3330.860 1711.920 ;
  LAYER metal2 ;
  RECT 3327.320 1710.800 3330.860 1711.920 ;
  LAYER metal1 ;
  RECT 3327.320 1710.800 3330.860 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3318.640 1710.800 3322.180 1711.920 ;
  LAYER metal4 ;
  RECT 3318.640 1710.800 3322.180 1711.920 ;
  LAYER metal3 ;
  RECT 3318.640 1710.800 3322.180 1711.920 ;
  LAYER metal2 ;
  RECT 3318.640 1710.800 3322.180 1711.920 ;
  LAYER metal1 ;
  RECT 3318.640 1710.800 3322.180 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3309.960 1710.800 3313.500 1711.920 ;
  LAYER metal4 ;
  RECT 3309.960 1710.800 3313.500 1711.920 ;
  LAYER metal3 ;
  RECT 3309.960 1710.800 3313.500 1711.920 ;
  LAYER metal2 ;
  RECT 3309.960 1710.800 3313.500 1711.920 ;
  LAYER metal1 ;
  RECT 3309.960 1710.800 3313.500 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3301.280 1710.800 3304.820 1711.920 ;
  LAYER metal4 ;
  RECT 3301.280 1710.800 3304.820 1711.920 ;
  LAYER metal3 ;
  RECT 3301.280 1710.800 3304.820 1711.920 ;
  LAYER metal2 ;
  RECT 3301.280 1710.800 3304.820 1711.920 ;
  LAYER metal1 ;
  RECT 3301.280 1710.800 3304.820 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3292.600 1710.800 3296.140 1711.920 ;
  LAYER metal4 ;
  RECT 3292.600 1710.800 3296.140 1711.920 ;
  LAYER metal3 ;
  RECT 3292.600 1710.800 3296.140 1711.920 ;
  LAYER metal2 ;
  RECT 3292.600 1710.800 3296.140 1711.920 ;
  LAYER metal1 ;
  RECT 3292.600 1710.800 3296.140 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3283.920 1710.800 3287.460 1711.920 ;
  LAYER metal4 ;
  RECT 3283.920 1710.800 3287.460 1711.920 ;
  LAYER metal3 ;
  RECT 3283.920 1710.800 3287.460 1711.920 ;
  LAYER metal2 ;
  RECT 3283.920 1710.800 3287.460 1711.920 ;
  LAYER metal1 ;
  RECT 3283.920 1710.800 3287.460 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3240.520 1710.800 3244.060 1711.920 ;
  LAYER metal4 ;
  RECT 3240.520 1710.800 3244.060 1711.920 ;
  LAYER metal3 ;
  RECT 3240.520 1710.800 3244.060 1711.920 ;
  LAYER metal2 ;
  RECT 3240.520 1710.800 3244.060 1711.920 ;
  LAYER metal1 ;
  RECT 3240.520 1710.800 3244.060 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3231.840 1710.800 3235.380 1711.920 ;
  LAYER metal4 ;
  RECT 3231.840 1710.800 3235.380 1711.920 ;
  LAYER metal3 ;
  RECT 3231.840 1710.800 3235.380 1711.920 ;
  LAYER metal2 ;
  RECT 3231.840 1710.800 3235.380 1711.920 ;
  LAYER metal1 ;
  RECT 3231.840 1710.800 3235.380 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3223.160 1710.800 3226.700 1711.920 ;
  LAYER metal4 ;
  RECT 3223.160 1710.800 3226.700 1711.920 ;
  LAYER metal3 ;
  RECT 3223.160 1710.800 3226.700 1711.920 ;
  LAYER metal2 ;
  RECT 3223.160 1710.800 3226.700 1711.920 ;
  LAYER metal1 ;
  RECT 3223.160 1710.800 3226.700 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3214.480 1710.800 3218.020 1711.920 ;
  LAYER metal4 ;
  RECT 3214.480 1710.800 3218.020 1711.920 ;
  LAYER metal3 ;
  RECT 3214.480 1710.800 3218.020 1711.920 ;
  LAYER metal2 ;
  RECT 3214.480 1710.800 3218.020 1711.920 ;
  LAYER metal1 ;
  RECT 3214.480 1710.800 3218.020 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3201.460 1710.800 3205.000 1711.920 ;
  LAYER metal4 ;
  RECT 3201.460 1710.800 3205.000 1711.920 ;
  LAYER metal3 ;
  RECT 3201.460 1710.800 3205.000 1711.920 ;
  LAYER metal2 ;
  RECT 3201.460 1710.800 3205.000 1711.920 ;
  LAYER metal1 ;
  RECT 3201.460 1710.800 3205.000 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3187.820 1710.800 3191.360 1711.920 ;
  LAYER metal4 ;
  RECT 3187.820 1710.800 3191.360 1711.920 ;
  LAYER metal3 ;
  RECT 3187.820 1710.800 3191.360 1711.920 ;
  LAYER metal2 ;
  RECT 3187.820 1710.800 3191.360 1711.920 ;
  LAYER metal1 ;
  RECT 3187.820 1710.800 3191.360 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3133.880 1710.800 3137.420 1711.920 ;
  LAYER metal4 ;
  RECT 3133.880 1710.800 3137.420 1711.920 ;
  LAYER metal3 ;
  RECT 3133.880 1710.800 3137.420 1711.920 ;
  LAYER metal2 ;
  RECT 3133.880 1710.800 3137.420 1711.920 ;
  LAYER metal1 ;
  RECT 3133.880 1710.800 3137.420 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3125.200 1710.800 3128.740 1711.920 ;
  LAYER metal4 ;
  RECT 3125.200 1710.800 3128.740 1711.920 ;
  LAYER metal3 ;
  RECT 3125.200 1710.800 3128.740 1711.920 ;
  LAYER metal2 ;
  RECT 3125.200 1710.800 3128.740 1711.920 ;
  LAYER metal1 ;
  RECT 3125.200 1710.800 3128.740 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3116.520 1710.800 3120.060 1711.920 ;
  LAYER metal4 ;
  RECT 3116.520 1710.800 3120.060 1711.920 ;
  LAYER metal3 ;
  RECT 3116.520 1710.800 3120.060 1711.920 ;
  LAYER metal2 ;
  RECT 3116.520 1710.800 3120.060 1711.920 ;
  LAYER metal1 ;
  RECT 3116.520 1710.800 3120.060 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3107.840 1710.800 3111.380 1711.920 ;
  LAYER metal4 ;
  RECT 3107.840 1710.800 3111.380 1711.920 ;
  LAYER metal3 ;
  RECT 3107.840 1710.800 3111.380 1711.920 ;
  LAYER metal2 ;
  RECT 3107.840 1710.800 3111.380 1711.920 ;
  LAYER metal1 ;
  RECT 3107.840 1710.800 3111.380 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3099.160 1710.800 3102.700 1711.920 ;
  LAYER metal4 ;
  RECT 3099.160 1710.800 3102.700 1711.920 ;
  LAYER metal3 ;
  RECT 3099.160 1710.800 3102.700 1711.920 ;
  LAYER metal2 ;
  RECT 3099.160 1710.800 3102.700 1711.920 ;
  LAYER metal1 ;
  RECT 3099.160 1710.800 3102.700 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3090.480 1710.800 3094.020 1711.920 ;
  LAYER metal4 ;
  RECT 3090.480 1710.800 3094.020 1711.920 ;
  LAYER metal3 ;
  RECT 3090.480 1710.800 3094.020 1711.920 ;
  LAYER metal2 ;
  RECT 3090.480 1710.800 3094.020 1711.920 ;
  LAYER metal1 ;
  RECT 3090.480 1710.800 3094.020 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3047.080 1710.800 3050.620 1711.920 ;
  LAYER metal4 ;
  RECT 3047.080 1710.800 3050.620 1711.920 ;
  LAYER metal3 ;
  RECT 3047.080 1710.800 3050.620 1711.920 ;
  LAYER metal2 ;
  RECT 3047.080 1710.800 3050.620 1711.920 ;
  LAYER metal1 ;
  RECT 3047.080 1710.800 3050.620 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3038.400 1710.800 3041.940 1711.920 ;
  LAYER metal4 ;
  RECT 3038.400 1710.800 3041.940 1711.920 ;
  LAYER metal3 ;
  RECT 3038.400 1710.800 3041.940 1711.920 ;
  LAYER metal2 ;
  RECT 3038.400 1710.800 3041.940 1711.920 ;
  LAYER metal1 ;
  RECT 3038.400 1710.800 3041.940 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3029.720 1710.800 3033.260 1711.920 ;
  LAYER metal4 ;
  RECT 3029.720 1710.800 3033.260 1711.920 ;
  LAYER metal3 ;
  RECT 3029.720 1710.800 3033.260 1711.920 ;
  LAYER metal2 ;
  RECT 3029.720 1710.800 3033.260 1711.920 ;
  LAYER metal1 ;
  RECT 3029.720 1710.800 3033.260 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3021.040 1710.800 3024.580 1711.920 ;
  LAYER metal4 ;
  RECT 3021.040 1710.800 3024.580 1711.920 ;
  LAYER metal3 ;
  RECT 3021.040 1710.800 3024.580 1711.920 ;
  LAYER metal2 ;
  RECT 3021.040 1710.800 3024.580 1711.920 ;
  LAYER metal1 ;
  RECT 3021.040 1710.800 3024.580 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3012.360 1710.800 3015.900 1711.920 ;
  LAYER metal4 ;
  RECT 3012.360 1710.800 3015.900 1711.920 ;
  LAYER metal3 ;
  RECT 3012.360 1710.800 3015.900 1711.920 ;
  LAYER metal2 ;
  RECT 3012.360 1710.800 3015.900 1711.920 ;
  LAYER metal1 ;
  RECT 3012.360 1710.800 3015.900 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3003.680 1710.800 3007.220 1711.920 ;
  LAYER metal4 ;
  RECT 3003.680 1710.800 3007.220 1711.920 ;
  LAYER metal3 ;
  RECT 3003.680 1710.800 3007.220 1711.920 ;
  LAYER metal2 ;
  RECT 3003.680 1710.800 3007.220 1711.920 ;
  LAYER metal1 ;
  RECT 3003.680 1710.800 3007.220 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2960.280 1710.800 2963.820 1711.920 ;
  LAYER metal4 ;
  RECT 2960.280 1710.800 2963.820 1711.920 ;
  LAYER metal3 ;
  RECT 2960.280 1710.800 2963.820 1711.920 ;
  LAYER metal2 ;
  RECT 2960.280 1710.800 2963.820 1711.920 ;
  LAYER metal1 ;
  RECT 2960.280 1710.800 2963.820 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2951.600 1710.800 2955.140 1711.920 ;
  LAYER metal4 ;
  RECT 2951.600 1710.800 2955.140 1711.920 ;
  LAYER metal3 ;
  RECT 2951.600 1710.800 2955.140 1711.920 ;
  LAYER metal2 ;
  RECT 2951.600 1710.800 2955.140 1711.920 ;
  LAYER metal1 ;
  RECT 2951.600 1710.800 2955.140 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2942.920 1710.800 2946.460 1711.920 ;
  LAYER metal4 ;
  RECT 2942.920 1710.800 2946.460 1711.920 ;
  LAYER metal3 ;
  RECT 2942.920 1710.800 2946.460 1711.920 ;
  LAYER metal2 ;
  RECT 2942.920 1710.800 2946.460 1711.920 ;
  LAYER metal1 ;
  RECT 2942.920 1710.800 2946.460 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2934.240 1710.800 2937.780 1711.920 ;
  LAYER metal4 ;
  RECT 2934.240 1710.800 2937.780 1711.920 ;
  LAYER metal3 ;
  RECT 2934.240 1710.800 2937.780 1711.920 ;
  LAYER metal2 ;
  RECT 2934.240 1710.800 2937.780 1711.920 ;
  LAYER metal1 ;
  RECT 2934.240 1710.800 2937.780 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2925.560 1710.800 2929.100 1711.920 ;
  LAYER metal4 ;
  RECT 2925.560 1710.800 2929.100 1711.920 ;
  LAYER metal3 ;
  RECT 2925.560 1710.800 2929.100 1711.920 ;
  LAYER metal2 ;
  RECT 2925.560 1710.800 2929.100 1711.920 ;
  LAYER metal1 ;
  RECT 2925.560 1710.800 2929.100 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2916.880 1710.800 2920.420 1711.920 ;
  LAYER metal4 ;
  RECT 2916.880 1710.800 2920.420 1711.920 ;
  LAYER metal3 ;
  RECT 2916.880 1710.800 2920.420 1711.920 ;
  LAYER metal2 ;
  RECT 2916.880 1710.800 2920.420 1711.920 ;
  LAYER metal1 ;
  RECT 2916.880 1710.800 2920.420 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2873.480 1710.800 2877.020 1711.920 ;
  LAYER metal4 ;
  RECT 2873.480 1710.800 2877.020 1711.920 ;
  LAYER metal3 ;
  RECT 2873.480 1710.800 2877.020 1711.920 ;
  LAYER metal2 ;
  RECT 2873.480 1710.800 2877.020 1711.920 ;
  LAYER metal1 ;
  RECT 2873.480 1710.800 2877.020 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2864.800 1710.800 2868.340 1711.920 ;
  LAYER metal4 ;
  RECT 2864.800 1710.800 2868.340 1711.920 ;
  LAYER metal3 ;
  RECT 2864.800 1710.800 2868.340 1711.920 ;
  LAYER metal2 ;
  RECT 2864.800 1710.800 2868.340 1711.920 ;
  LAYER metal1 ;
  RECT 2864.800 1710.800 2868.340 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2856.120 1710.800 2859.660 1711.920 ;
  LAYER metal4 ;
  RECT 2856.120 1710.800 2859.660 1711.920 ;
  LAYER metal3 ;
  RECT 2856.120 1710.800 2859.660 1711.920 ;
  LAYER metal2 ;
  RECT 2856.120 1710.800 2859.660 1711.920 ;
  LAYER metal1 ;
  RECT 2856.120 1710.800 2859.660 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2847.440 1710.800 2850.980 1711.920 ;
  LAYER metal4 ;
  RECT 2847.440 1710.800 2850.980 1711.920 ;
  LAYER metal3 ;
  RECT 2847.440 1710.800 2850.980 1711.920 ;
  LAYER metal2 ;
  RECT 2847.440 1710.800 2850.980 1711.920 ;
  LAYER metal1 ;
  RECT 2847.440 1710.800 2850.980 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2838.760 1710.800 2842.300 1711.920 ;
  LAYER metal4 ;
  RECT 2838.760 1710.800 2842.300 1711.920 ;
  LAYER metal3 ;
  RECT 2838.760 1710.800 2842.300 1711.920 ;
  LAYER metal2 ;
  RECT 2838.760 1710.800 2842.300 1711.920 ;
  LAYER metal1 ;
  RECT 2838.760 1710.800 2842.300 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2830.080 1710.800 2833.620 1711.920 ;
  LAYER metal4 ;
  RECT 2830.080 1710.800 2833.620 1711.920 ;
  LAYER metal3 ;
  RECT 2830.080 1710.800 2833.620 1711.920 ;
  LAYER metal2 ;
  RECT 2830.080 1710.800 2833.620 1711.920 ;
  LAYER metal1 ;
  RECT 2830.080 1710.800 2833.620 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2786.680 1710.800 2790.220 1711.920 ;
  LAYER metal4 ;
  RECT 2786.680 1710.800 2790.220 1711.920 ;
  LAYER metal3 ;
  RECT 2786.680 1710.800 2790.220 1711.920 ;
  LAYER metal2 ;
  RECT 2786.680 1710.800 2790.220 1711.920 ;
  LAYER metal1 ;
  RECT 2786.680 1710.800 2790.220 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2773.660 1710.800 2777.200 1711.920 ;
  LAYER metal4 ;
  RECT 2773.660 1710.800 2777.200 1711.920 ;
  LAYER metal3 ;
  RECT 2773.660 1710.800 2777.200 1711.920 ;
  LAYER metal2 ;
  RECT 2773.660 1710.800 2777.200 1711.920 ;
  LAYER metal1 ;
  RECT 2773.660 1710.800 2777.200 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2760.020 1710.800 2763.560 1711.920 ;
  LAYER metal4 ;
  RECT 2760.020 1710.800 2763.560 1711.920 ;
  LAYER metal3 ;
  RECT 2760.020 1710.800 2763.560 1711.920 ;
  LAYER metal2 ;
  RECT 2760.020 1710.800 2763.560 1711.920 ;
  LAYER metal1 ;
  RECT 2760.020 1710.800 2763.560 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2746.380 1710.800 2749.920 1711.920 ;
  LAYER metal4 ;
  RECT 2746.380 1710.800 2749.920 1711.920 ;
  LAYER metal3 ;
  RECT 2746.380 1710.800 2749.920 1711.920 ;
  LAYER metal2 ;
  RECT 2746.380 1710.800 2749.920 1711.920 ;
  LAYER metal1 ;
  RECT 2746.380 1710.800 2749.920 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2732.120 1710.800 2735.660 1711.920 ;
  LAYER metal4 ;
  RECT 2732.120 1710.800 2735.660 1711.920 ;
  LAYER metal3 ;
  RECT 2732.120 1710.800 2735.660 1711.920 ;
  LAYER metal2 ;
  RECT 2732.120 1710.800 2735.660 1711.920 ;
  LAYER metal1 ;
  RECT 2732.120 1710.800 2735.660 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2723.440 1710.800 2726.980 1711.920 ;
  LAYER metal4 ;
  RECT 2723.440 1710.800 2726.980 1711.920 ;
  LAYER metal3 ;
  RECT 2723.440 1710.800 2726.980 1711.920 ;
  LAYER metal2 ;
  RECT 2723.440 1710.800 2726.980 1711.920 ;
  LAYER metal1 ;
  RECT 2723.440 1710.800 2726.980 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2680.040 1710.800 2683.580 1711.920 ;
  LAYER metal4 ;
  RECT 2680.040 1710.800 2683.580 1711.920 ;
  LAYER metal3 ;
  RECT 2680.040 1710.800 2683.580 1711.920 ;
  LAYER metal2 ;
  RECT 2680.040 1710.800 2683.580 1711.920 ;
  LAYER metal1 ;
  RECT 2680.040 1710.800 2683.580 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2671.360 1710.800 2674.900 1711.920 ;
  LAYER metal4 ;
  RECT 2671.360 1710.800 2674.900 1711.920 ;
  LAYER metal3 ;
  RECT 2671.360 1710.800 2674.900 1711.920 ;
  LAYER metal2 ;
  RECT 2671.360 1710.800 2674.900 1711.920 ;
  LAYER metal1 ;
  RECT 2671.360 1710.800 2674.900 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2662.680 1710.800 2666.220 1711.920 ;
  LAYER metal4 ;
  RECT 2662.680 1710.800 2666.220 1711.920 ;
  LAYER metal3 ;
  RECT 2662.680 1710.800 2666.220 1711.920 ;
  LAYER metal2 ;
  RECT 2662.680 1710.800 2666.220 1711.920 ;
  LAYER metal1 ;
  RECT 2662.680 1710.800 2666.220 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2654.000 1710.800 2657.540 1711.920 ;
  LAYER metal4 ;
  RECT 2654.000 1710.800 2657.540 1711.920 ;
  LAYER metal3 ;
  RECT 2654.000 1710.800 2657.540 1711.920 ;
  LAYER metal2 ;
  RECT 2654.000 1710.800 2657.540 1711.920 ;
  LAYER metal1 ;
  RECT 2654.000 1710.800 2657.540 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2645.320 1710.800 2648.860 1711.920 ;
  LAYER metal4 ;
  RECT 2645.320 1710.800 2648.860 1711.920 ;
  LAYER metal3 ;
  RECT 2645.320 1710.800 2648.860 1711.920 ;
  LAYER metal2 ;
  RECT 2645.320 1710.800 2648.860 1711.920 ;
  LAYER metal1 ;
  RECT 2645.320 1710.800 2648.860 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2636.640 1710.800 2640.180 1711.920 ;
  LAYER metal4 ;
  RECT 2636.640 1710.800 2640.180 1711.920 ;
  LAYER metal3 ;
  RECT 2636.640 1710.800 2640.180 1711.920 ;
  LAYER metal2 ;
  RECT 2636.640 1710.800 2640.180 1711.920 ;
  LAYER metal1 ;
  RECT 2636.640 1710.800 2640.180 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2593.240 1710.800 2596.780 1711.920 ;
  LAYER metal4 ;
  RECT 2593.240 1710.800 2596.780 1711.920 ;
  LAYER metal3 ;
  RECT 2593.240 1710.800 2596.780 1711.920 ;
  LAYER metal2 ;
  RECT 2593.240 1710.800 2596.780 1711.920 ;
  LAYER metal1 ;
  RECT 2593.240 1710.800 2596.780 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2584.560 1710.800 2588.100 1711.920 ;
  LAYER metal4 ;
  RECT 2584.560 1710.800 2588.100 1711.920 ;
  LAYER metal3 ;
  RECT 2584.560 1710.800 2588.100 1711.920 ;
  LAYER metal2 ;
  RECT 2584.560 1710.800 2588.100 1711.920 ;
  LAYER metal1 ;
  RECT 2584.560 1710.800 2588.100 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2575.880 1710.800 2579.420 1711.920 ;
  LAYER metal4 ;
  RECT 2575.880 1710.800 2579.420 1711.920 ;
  LAYER metal3 ;
  RECT 2575.880 1710.800 2579.420 1711.920 ;
  LAYER metal2 ;
  RECT 2575.880 1710.800 2579.420 1711.920 ;
  LAYER metal1 ;
  RECT 2575.880 1710.800 2579.420 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2567.200 1710.800 2570.740 1711.920 ;
  LAYER metal4 ;
  RECT 2567.200 1710.800 2570.740 1711.920 ;
  LAYER metal3 ;
  RECT 2567.200 1710.800 2570.740 1711.920 ;
  LAYER metal2 ;
  RECT 2567.200 1710.800 2570.740 1711.920 ;
  LAYER metal1 ;
  RECT 2567.200 1710.800 2570.740 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2558.520 1710.800 2562.060 1711.920 ;
  LAYER metal4 ;
  RECT 2558.520 1710.800 2562.060 1711.920 ;
  LAYER metal3 ;
  RECT 2558.520 1710.800 2562.060 1711.920 ;
  LAYER metal2 ;
  RECT 2558.520 1710.800 2562.060 1711.920 ;
  LAYER metal1 ;
  RECT 2558.520 1710.800 2562.060 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2549.840 1710.800 2553.380 1711.920 ;
  LAYER metal4 ;
  RECT 2549.840 1710.800 2553.380 1711.920 ;
  LAYER metal3 ;
  RECT 2549.840 1710.800 2553.380 1711.920 ;
  LAYER metal2 ;
  RECT 2549.840 1710.800 2553.380 1711.920 ;
  LAYER metal1 ;
  RECT 2549.840 1710.800 2553.380 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2506.440 1710.800 2509.980 1711.920 ;
  LAYER metal4 ;
  RECT 2506.440 1710.800 2509.980 1711.920 ;
  LAYER metal3 ;
  RECT 2506.440 1710.800 2509.980 1711.920 ;
  LAYER metal2 ;
  RECT 2506.440 1710.800 2509.980 1711.920 ;
  LAYER metal1 ;
  RECT 2506.440 1710.800 2509.980 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2497.760 1710.800 2501.300 1711.920 ;
  LAYER metal4 ;
  RECT 2497.760 1710.800 2501.300 1711.920 ;
  LAYER metal3 ;
  RECT 2497.760 1710.800 2501.300 1711.920 ;
  LAYER metal2 ;
  RECT 2497.760 1710.800 2501.300 1711.920 ;
  LAYER metal1 ;
  RECT 2497.760 1710.800 2501.300 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2489.080 1710.800 2492.620 1711.920 ;
  LAYER metal4 ;
  RECT 2489.080 1710.800 2492.620 1711.920 ;
  LAYER metal3 ;
  RECT 2489.080 1710.800 2492.620 1711.920 ;
  LAYER metal2 ;
  RECT 2489.080 1710.800 2492.620 1711.920 ;
  LAYER metal1 ;
  RECT 2489.080 1710.800 2492.620 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2480.400 1710.800 2483.940 1711.920 ;
  LAYER metal4 ;
  RECT 2480.400 1710.800 2483.940 1711.920 ;
  LAYER metal3 ;
  RECT 2480.400 1710.800 2483.940 1711.920 ;
  LAYER metal2 ;
  RECT 2480.400 1710.800 2483.940 1711.920 ;
  LAYER metal1 ;
  RECT 2480.400 1710.800 2483.940 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2471.720 1710.800 2475.260 1711.920 ;
  LAYER metal4 ;
  RECT 2471.720 1710.800 2475.260 1711.920 ;
  LAYER metal3 ;
  RECT 2471.720 1710.800 2475.260 1711.920 ;
  LAYER metal2 ;
  RECT 2471.720 1710.800 2475.260 1711.920 ;
  LAYER metal1 ;
  RECT 2471.720 1710.800 2475.260 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2463.040 1710.800 2466.580 1711.920 ;
  LAYER metal4 ;
  RECT 2463.040 1710.800 2466.580 1711.920 ;
  LAYER metal3 ;
  RECT 2463.040 1710.800 2466.580 1711.920 ;
  LAYER metal2 ;
  RECT 2463.040 1710.800 2466.580 1711.920 ;
  LAYER metal1 ;
  RECT 2463.040 1710.800 2466.580 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2419.640 1710.800 2423.180 1711.920 ;
  LAYER metal4 ;
  RECT 2419.640 1710.800 2423.180 1711.920 ;
  LAYER metal3 ;
  RECT 2419.640 1710.800 2423.180 1711.920 ;
  LAYER metal2 ;
  RECT 2419.640 1710.800 2423.180 1711.920 ;
  LAYER metal1 ;
  RECT 2419.640 1710.800 2423.180 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2410.960 1710.800 2414.500 1711.920 ;
  LAYER metal4 ;
  RECT 2410.960 1710.800 2414.500 1711.920 ;
  LAYER metal3 ;
  RECT 2410.960 1710.800 2414.500 1711.920 ;
  LAYER metal2 ;
  RECT 2410.960 1710.800 2414.500 1711.920 ;
  LAYER metal1 ;
  RECT 2410.960 1710.800 2414.500 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2402.280 1710.800 2405.820 1711.920 ;
  LAYER metal4 ;
  RECT 2402.280 1710.800 2405.820 1711.920 ;
  LAYER metal3 ;
  RECT 2402.280 1710.800 2405.820 1711.920 ;
  LAYER metal2 ;
  RECT 2402.280 1710.800 2405.820 1711.920 ;
  LAYER metal1 ;
  RECT 2402.280 1710.800 2405.820 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2393.600 1710.800 2397.140 1711.920 ;
  LAYER metal4 ;
  RECT 2393.600 1710.800 2397.140 1711.920 ;
  LAYER metal3 ;
  RECT 2393.600 1710.800 2397.140 1711.920 ;
  LAYER metal2 ;
  RECT 2393.600 1710.800 2397.140 1711.920 ;
  LAYER metal1 ;
  RECT 2393.600 1710.800 2397.140 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2384.920 1710.800 2388.460 1711.920 ;
  LAYER metal4 ;
  RECT 2384.920 1710.800 2388.460 1711.920 ;
  LAYER metal3 ;
  RECT 2384.920 1710.800 2388.460 1711.920 ;
  LAYER metal2 ;
  RECT 2384.920 1710.800 2388.460 1711.920 ;
  LAYER metal1 ;
  RECT 2384.920 1710.800 2388.460 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2376.240 1710.800 2379.780 1711.920 ;
  LAYER metal4 ;
  RECT 2376.240 1710.800 2379.780 1711.920 ;
  LAYER metal3 ;
  RECT 2376.240 1710.800 2379.780 1711.920 ;
  LAYER metal2 ;
  RECT 2376.240 1710.800 2379.780 1711.920 ;
  LAYER metal1 ;
  RECT 2376.240 1710.800 2379.780 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2323.540 1710.800 2327.080 1711.920 ;
  LAYER metal4 ;
  RECT 2323.540 1710.800 2327.080 1711.920 ;
  LAYER metal3 ;
  RECT 2323.540 1710.800 2327.080 1711.920 ;
  LAYER metal2 ;
  RECT 2323.540 1710.800 2327.080 1711.920 ;
  LAYER metal1 ;
  RECT 2323.540 1710.800 2327.080 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2309.900 1710.800 2313.440 1711.920 ;
  LAYER metal4 ;
  RECT 2309.900 1710.800 2313.440 1711.920 ;
  LAYER metal3 ;
  RECT 2309.900 1710.800 2313.440 1711.920 ;
  LAYER metal2 ;
  RECT 2309.900 1710.800 2313.440 1711.920 ;
  LAYER metal1 ;
  RECT 2309.900 1710.800 2313.440 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2295.640 1710.800 2299.180 1711.920 ;
  LAYER metal4 ;
  RECT 2295.640 1710.800 2299.180 1711.920 ;
  LAYER metal3 ;
  RECT 2295.640 1710.800 2299.180 1711.920 ;
  LAYER metal2 ;
  RECT 2295.640 1710.800 2299.180 1711.920 ;
  LAYER metal1 ;
  RECT 2295.640 1710.800 2299.180 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2286.960 1710.800 2290.500 1711.920 ;
  LAYER metal4 ;
  RECT 2286.960 1710.800 2290.500 1711.920 ;
  LAYER metal3 ;
  RECT 2286.960 1710.800 2290.500 1711.920 ;
  LAYER metal2 ;
  RECT 2286.960 1710.800 2290.500 1711.920 ;
  LAYER metal1 ;
  RECT 2286.960 1710.800 2290.500 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2278.280 1710.800 2281.820 1711.920 ;
  LAYER metal4 ;
  RECT 2278.280 1710.800 2281.820 1711.920 ;
  LAYER metal3 ;
  RECT 2278.280 1710.800 2281.820 1711.920 ;
  LAYER metal2 ;
  RECT 2278.280 1710.800 2281.820 1711.920 ;
  LAYER metal1 ;
  RECT 2278.280 1710.800 2281.820 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2269.600 1710.800 2273.140 1711.920 ;
  LAYER metal4 ;
  RECT 2269.600 1710.800 2273.140 1711.920 ;
  LAYER metal3 ;
  RECT 2269.600 1710.800 2273.140 1711.920 ;
  LAYER metal2 ;
  RECT 2269.600 1710.800 2273.140 1711.920 ;
  LAYER metal1 ;
  RECT 2269.600 1710.800 2273.140 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2226.200 1710.800 2229.740 1711.920 ;
  LAYER metal4 ;
  RECT 2226.200 1710.800 2229.740 1711.920 ;
  LAYER metal3 ;
  RECT 2226.200 1710.800 2229.740 1711.920 ;
  LAYER metal2 ;
  RECT 2226.200 1710.800 2229.740 1711.920 ;
  LAYER metal1 ;
  RECT 2226.200 1710.800 2229.740 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2217.520 1710.800 2221.060 1711.920 ;
  LAYER metal4 ;
  RECT 2217.520 1710.800 2221.060 1711.920 ;
  LAYER metal3 ;
  RECT 2217.520 1710.800 2221.060 1711.920 ;
  LAYER metal2 ;
  RECT 2217.520 1710.800 2221.060 1711.920 ;
  LAYER metal1 ;
  RECT 2217.520 1710.800 2221.060 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2208.840 1710.800 2212.380 1711.920 ;
  LAYER metal4 ;
  RECT 2208.840 1710.800 2212.380 1711.920 ;
  LAYER metal3 ;
  RECT 2208.840 1710.800 2212.380 1711.920 ;
  LAYER metal2 ;
  RECT 2208.840 1710.800 2212.380 1711.920 ;
  LAYER metal1 ;
  RECT 2208.840 1710.800 2212.380 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2200.160 1710.800 2203.700 1711.920 ;
  LAYER metal4 ;
  RECT 2200.160 1710.800 2203.700 1711.920 ;
  LAYER metal3 ;
  RECT 2200.160 1710.800 2203.700 1711.920 ;
  LAYER metal2 ;
  RECT 2200.160 1710.800 2203.700 1711.920 ;
  LAYER metal1 ;
  RECT 2200.160 1710.800 2203.700 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2191.480 1710.800 2195.020 1711.920 ;
  LAYER metal4 ;
  RECT 2191.480 1710.800 2195.020 1711.920 ;
  LAYER metal3 ;
  RECT 2191.480 1710.800 2195.020 1711.920 ;
  LAYER metal2 ;
  RECT 2191.480 1710.800 2195.020 1711.920 ;
  LAYER metal1 ;
  RECT 2191.480 1710.800 2195.020 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2182.800 1710.800 2186.340 1711.920 ;
  LAYER metal4 ;
  RECT 2182.800 1710.800 2186.340 1711.920 ;
  LAYER metal3 ;
  RECT 2182.800 1710.800 2186.340 1711.920 ;
  LAYER metal2 ;
  RECT 2182.800 1710.800 2186.340 1711.920 ;
  LAYER metal1 ;
  RECT 2182.800 1710.800 2186.340 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2139.400 1710.800 2142.940 1711.920 ;
  LAYER metal4 ;
  RECT 2139.400 1710.800 2142.940 1711.920 ;
  LAYER metal3 ;
  RECT 2139.400 1710.800 2142.940 1711.920 ;
  LAYER metal2 ;
  RECT 2139.400 1710.800 2142.940 1711.920 ;
  LAYER metal1 ;
  RECT 2139.400 1710.800 2142.940 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2130.720 1710.800 2134.260 1711.920 ;
  LAYER metal4 ;
  RECT 2130.720 1710.800 2134.260 1711.920 ;
  LAYER metal3 ;
  RECT 2130.720 1710.800 2134.260 1711.920 ;
  LAYER metal2 ;
  RECT 2130.720 1710.800 2134.260 1711.920 ;
  LAYER metal1 ;
  RECT 2130.720 1710.800 2134.260 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2122.040 1710.800 2125.580 1711.920 ;
  LAYER metal4 ;
  RECT 2122.040 1710.800 2125.580 1711.920 ;
  LAYER metal3 ;
  RECT 2122.040 1710.800 2125.580 1711.920 ;
  LAYER metal2 ;
  RECT 2122.040 1710.800 2125.580 1711.920 ;
  LAYER metal1 ;
  RECT 2122.040 1710.800 2125.580 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2113.360 1710.800 2116.900 1711.920 ;
  LAYER metal4 ;
  RECT 2113.360 1710.800 2116.900 1711.920 ;
  LAYER metal3 ;
  RECT 2113.360 1710.800 2116.900 1711.920 ;
  LAYER metal2 ;
  RECT 2113.360 1710.800 2116.900 1711.920 ;
  LAYER metal1 ;
  RECT 2113.360 1710.800 2116.900 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2104.680 1710.800 2108.220 1711.920 ;
  LAYER metal4 ;
  RECT 2104.680 1710.800 2108.220 1711.920 ;
  LAYER metal3 ;
  RECT 2104.680 1710.800 2108.220 1711.920 ;
  LAYER metal2 ;
  RECT 2104.680 1710.800 2108.220 1711.920 ;
  LAYER metal1 ;
  RECT 2104.680 1710.800 2108.220 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2096.000 1710.800 2099.540 1711.920 ;
  LAYER metal4 ;
  RECT 2096.000 1710.800 2099.540 1711.920 ;
  LAYER metal3 ;
  RECT 2096.000 1710.800 2099.540 1711.920 ;
  LAYER metal2 ;
  RECT 2096.000 1710.800 2099.540 1711.920 ;
  LAYER metal1 ;
  RECT 2096.000 1710.800 2099.540 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2052.600 1710.800 2056.140 1711.920 ;
  LAYER metal4 ;
  RECT 2052.600 1710.800 2056.140 1711.920 ;
  LAYER metal3 ;
  RECT 2052.600 1710.800 2056.140 1711.920 ;
  LAYER metal2 ;
  RECT 2052.600 1710.800 2056.140 1711.920 ;
  LAYER metal1 ;
  RECT 2052.600 1710.800 2056.140 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2043.920 1710.800 2047.460 1711.920 ;
  LAYER metal4 ;
  RECT 2043.920 1710.800 2047.460 1711.920 ;
  LAYER metal3 ;
  RECT 2043.920 1710.800 2047.460 1711.920 ;
  LAYER metal2 ;
  RECT 2043.920 1710.800 2047.460 1711.920 ;
  LAYER metal1 ;
  RECT 2043.920 1710.800 2047.460 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2035.240 1710.800 2038.780 1711.920 ;
  LAYER metal4 ;
  RECT 2035.240 1710.800 2038.780 1711.920 ;
  LAYER metal3 ;
  RECT 2035.240 1710.800 2038.780 1711.920 ;
  LAYER metal2 ;
  RECT 2035.240 1710.800 2038.780 1711.920 ;
  LAYER metal1 ;
  RECT 2035.240 1710.800 2038.780 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2026.560 1710.800 2030.100 1711.920 ;
  LAYER metal4 ;
  RECT 2026.560 1710.800 2030.100 1711.920 ;
  LAYER metal3 ;
  RECT 2026.560 1710.800 2030.100 1711.920 ;
  LAYER metal2 ;
  RECT 2026.560 1710.800 2030.100 1711.920 ;
  LAYER metal1 ;
  RECT 2026.560 1710.800 2030.100 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2017.880 1710.800 2021.420 1711.920 ;
  LAYER metal4 ;
  RECT 2017.880 1710.800 2021.420 1711.920 ;
  LAYER metal3 ;
  RECT 2017.880 1710.800 2021.420 1711.920 ;
  LAYER metal2 ;
  RECT 2017.880 1710.800 2021.420 1711.920 ;
  LAYER metal1 ;
  RECT 2017.880 1710.800 2021.420 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2009.200 1710.800 2012.740 1711.920 ;
  LAYER metal4 ;
  RECT 2009.200 1710.800 2012.740 1711.920 ;
  LAYER metal3 ;
  RECT 2009.200 1710.800 2012.740 1711.920 ;
  LAYER metal2 ;
  RECT 2009.200 1710.800 2012.740 1711.920 ;
  LAYER metal1 ;
  RECT 2009.200 1710.800 2012.740 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1965.800 1710.800 1969.340 1711.920 ;
  LAYER metal4 ;
  RECT 1965.800 1710.800 1969.340 1711.920 ;
  LAYER metal3 ;
  RECT 1965.800 1710.800 1969.340 1711.920 ;
  LAYER metal2 ;
  RECT 1965.800 1710.800 1969.340 1711.920 ;
  LAYER metal1 ;
  RECT 1965.800 1710.800 1969.340 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1957.120 1710.800 1960.660 1711.920 ;
  LAYER metal4 ;
  RECT 1957.120 1710.800 1960.660 1711.920 ;
  LAYER metal3 ;
  RECT 1957.120 1710.800 1960.660 1711.920 ;
  LAYER metal2 ;
  RECT 1957.120 1710.800 1960.660 1711.920 ;
  LAYER metal1 ;
  RECT 1957.120 1710.800 1960.660 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1948.440 1710.800 1951.980 1711.920 ;
  LAYER metal4 ;
  RECT 1948.440 1710.800 1951.980 1711.920 ;
  LAYER metal3 ;
  RECT 1948.440 1710.800 1951.980 1711.920 ;
  LAYER metal2 ;
  RECT 1948.440 1710.800 1951.980 1711.920 ;
  LAYER metal1 ;
  RECT 1948.440 1710.800 1951.980 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1939.760 1710.800 1943.300 1711.920 ;
  LAYER metal4 ;
  RECT 1939.760 1710.800 1943.300 1711.920 ;
  LAYER metal3 ;
  RECT 1939.760 1710.800 1943.300 1711.920 ;
  LAYER metal2 ;
  RECT 1939.760 1710.800 1943.300 1711.920 ;
  LAYER metal1 ;
  RECT 1939.760 1710.800 1943.300 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1931.080 1710.800 1934.620 1711.920 ;
  LAYER metal4 ;
  RECT 1931.080 1710.800 1934.620 1711.920 ;
  LAYER metal3 ;
  RECT 1931.080 1710.800 1934.620 1711.920 ;
  LAYER metal2 ;
  RECT 1931.080 1710.800 1934.620 1711.920 ;
  LAYER metal1 ;
  RECT 1931.080 1710.800 1934.620 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1922.400 1710.800 1925.940 1711.920 ;
  LAYER metal4 ;
  RECT 1922.400 1710.800 1925.940 1711.920 ;
  LAYER metal3 ;
  RECT 1922.400 1710.800 1925.940 1711.920 ;
  LAYER metal2 ;
  RECT 1922.400 1710.800 1925.940 1711.920 ;
  LAYER metal1 ;
  RECT 1922.400 1710.800 1925.940 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1859.160 1710.800 1862.700 1711.920 ;
  LAYER metal4 ;
  RECT 1859.160 1710.800 1862.700 1711.920 ;
  LAYER metal3 ;
  RECT 1859.160 1710.800 1862.700 1711.920 ;
  LAYER metal2 ;
  RECT 1859.160 1710.800 1862.700 1711.920 ;
  LAYER metal1 ;
  RECT 1859.160 1710.800 1862.700 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1850.480 1710.800 1854.020 1711.920 ;
  LAYER metal4 ;
  RECT 1850.480 1710.800 1854.020 1711.920 ;
  LAYER metal3 ;
  RECT 1850.480 1710.800 1854.020 1711.920 ;
  LAYER metal2 ;
  RECT 1850.480 1710.800 1854.020 1711.920 ;
  LAYER metal1 ;
  RECT 1850.480 1710.800 1854.020 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1793.440 1710.800 1796.980 1711.920 ;
  LAYER metal4 ;
  RECT 1793.440 1710.800 1796.980 1711.920 ;
  LAYER metal3 ;
  RECT 1793.440 1710.800 1796.980 1711.920 ;
  LAYER metal2 ;
  RECT 1793.440 1710.800 1796.980 1711.920 ;
  LAYER metal1 ;
  RECT 1793.440 1710.800 1796.980 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1768.640 1710.800 1772.180 1711.920 ;
  LAYER metal4 ;
  RECT 1768.640 1710.800 1772.180 1711.920 ;
  LAYER metal3 ;
  RECT 1768.640 1710.800 1772.180 1711.920 ;
  LAYER metal2 ;
  RECT 1768.640 1710.800 1772.180 1711.920 ;
  LAYER metal1 ;
  RECT 1768.640 1710.800 1772.180 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1742.600 1710.800 1746.140 1711.920 ;
  LAYER metal4 ;
  RECT 1742.600 1710.800 1746.140 1711.920 ;
  LAYER metal3 ;
  RECT 1742.600 1710.800 1746.140 1711.920 ;
  LAYER metal2 ;
  RECT 1742.600 1710.800 1746.140 1711.920 ;
  LAYER metal1 ;
  RECT 1742.600 1710.800 1746.140 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1733.920 1710.800 1737.460 1711.920 ;
  LAYER metal4 ;
  RECT 1733.920 1710.800 1737.460 1711.920 ;
  LAYER metal3 ;
  RECT 1733.920 1710.800 1737.460 1711.920 ;
  LAYER metal2 ;
  RECT 1733.920 1710.800 1737.460 1711.920 ;
  LAYER metal1 ;
  RECT 1733.920 1710.800 1737.460 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1690.520 1710.800 1694.060 1711.920 ;
  LAYER metal4 ;
  RECT 1690.520 1710.800 1694.060 1711.920 ;
  LAYER metal3 ;
  RECT 1690.520 1710.800 1694.060 1711.920 ;
  LAYER metal2 ;
  RECT 1690.520 1710.800 1694.060 1711.920 ;
  LAYER metal1 ;
  RECT 1690.520 1710.800 1694.060 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1681.840 1710.800 1685.380 1711.920 ;
  LAYER metal4 ;
  RECT 1681.840 1710.800 1685.380 1711.920 ;
  LAYER metal3 ;
  RECT 1681.840 1710.800 1685.380 1711.920 ;
  LAYER metal2 ;
  RECT 1681.840 1710.800 1685.380 1711.920 ;
  LAYER metal1 ;
  RECT 1681.840 1710.800 1685.380 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1673.160 1710.800 1676.700 1711.920 ;
  LAYER metal4 ;
  RECT 1673.160 1710.800 1676.700 1711.920 ;
  LAYER metal3 ;
  RECT 1673.160 1710.800 1676.700 1711.920 ;
  LAYER metal2 ;
  RECT 1673.160 1710.800 1676.700 1711.920 ;
  LAYER metal1 ;
  RECT 1673.160 1710.800 1676.700 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1664.480 1710.800 1668.020 1711.920 ;
  LAYER metal4 ;
  RECT 1664.480 1710.800 1668.020 1711.920 ;
  LAYER metal3 ;
  RECT 1664.480 1710.800 1668.020 1711.920 ;
  LAYER metal2 ;
  RECT 1664.480 1710.800 1668.020 1711.920 ;
  LAYER metal1 ;
  RECT 1664.480 1710.800 1668.020 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1655.800 1710.800 1659.340 1711.920 ;
  LAYER metal4 ;
  RECT 1655.800 1710.800 1659.340 1711.920 ;
  LAYER metal3 ;
  RECT 1655.800 1710.800 1659.340 1711.920 ;
  LAYER metal2 ;
  RECT 1655.800 1710.800 1659.340 1711.920 ;
  LAYER metal1 ;
  RECT 1655.800 1710.800 1659.340 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1647.120 1710.800 1650.660 1711.920 ;
  LAYER metal4 ;
  RECT 1647.120 1710.800 1650.660 1711.920 ;
  LAYER metal3 ;
  RECT 1647.120 1710.800 1650.660 1711.920 ;
  LAYER metal2 ;
  RECT 1647.120 1710.800 1650.660 1711.920 ;
  LAYER metal1 ;
  RECT 1647.120 1710.800 1650.660 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1603.720 1710.800 1607.260 1711.920 ;
  LAYER metal4 ;
  RECT 1603.720 1710.800 1607.260 1711.920 ;
  LAYER metal3 ;
  RECT 1603.720 1710.800 1607.260 1711.920 ;
  LAYER metal2 ;
  RECT 1603.720 1710.800 1607.260 1711.920 ;
  LAYER metal1 ;
  RECT 1603.720 1710.800 1607.260 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1595.040 1710.800 1598.580 1711.920 ;
  LAYER metal4 ;
  RECT 1595.040 1710.800 1598.580 1711.920 ;
  LAYER metal3 ;
  RECT 1595.040 1710.800 1598.580 1711.920 ;
  LAYER metal2 ;
  RECT 1595.040 1710.800 1598.580 1711.920 ;
  LAYER metal1 ;
  RECT 1595.040 1710.800 1598.580 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1586.360 1710.800 1589.900 1711.920 ;
  LAYER metal4 ;
  RECT 1586.360 1710.800 1589.900 1711.920 ;
  LAYER metal3 ;
  RECT 1586.360 1710.800 1589.900 1711.920 ;
  LAYER metal2 ;
  RECT 1586.360 1710.800 1589.900 1711.920 ;
  LAYER metal1 ;
  RECT 1586.360 1710.800 1589.900 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1577.680 1710.800 1581.220 1711.920 ;
  LAYER metal4 ;
  RECT 1577.680 1710.800 1581.220 1711.920 ;
  LAYER metal3 ;
  RECT 1577.680 1710.800 1581.220 1711.920 ;
  LAYER metal2 ;
  RECT 1577.680 1710.800 1581.220 1711.920 ;
  LAYER metal1 ;
  RECT 1577.680 1710.800 1581.220 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1569.000 1710.800 1572.540 1711.920 ;
  LAYER metal4 ;
  RECT 1569.000 1710.800 1572.540 1711.920 ;
  LAYER metal3 ;
  RECT 1569.000 1710.800 1572.540 1711.920 ;
  LAYER metal2 ;
  RECT 1569.000 1710.800 1572.540 1711.920 ;
  LAYER metal1 ;
  RECT 1569.000 1710.800 1572.540 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1560.320 1710.800 1563.860 1711.920 ;
  LAYER metal4 ;
  RECT 1560.320 1710.800 1563.860 1711.920 ;
  LAYER metal3 ;
  RECT 1560.320 1710.800 1563.860 1711.920 ;
  LAYER metal2 ;
  RECT 1560.320 1710.800 1563.860 1711.920 ;
  LAYER metal1 ;
  RECT 1560.320 1710.800 1563.860 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1516.920 1710.800 1520.460 1711.920 ;
  LAYER metal4 ;
  RECT 1516.920 1710.800 1520.460 1711.920 ;
  LAYER metal3 ;
  RECT 1516.920 1710.800 1520.460 1711.920 ;
  LAYER metal2 ;
  RECT 1516.920 1710.800 1520.460 1711.920 ;
  LAYER metal1 ;
  RECT 1516.920 1710.800 1520.460 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1508.240 1710.800 1511.780 1711.920 ;
  LAYER metal4 ;
  RECT 1508.240 1710.800 1511.780 1711.920 ;
  LAYER metal3 ;
  RECT 1508.240 1710.800 1511.780 1711.920 ;
  LAYER metal2 ;
  RECT 1508.240 1710.800 1511.780 1711.920 ;
  LAYER metal1 ;
  RECT 1508.240 1710.800 1511.780 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1499.560 1710.800 1503.100 1711.920 ;
  LAYER metal4 ;
  RECT 1499.560 1710.800 1503.100 1711.920 ;
  LAYER metal3 ;
  RECT 1499.560 1710.800 1503.100 1711.920 ;
  LAYER metal2 ;
  RECT 1499.560 1710.800 1503.100 1711.920 ;
  LAYER metal1 ;
  RECT 1499.560 1710.800 1503.100 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1490.880 1710.800 1494.420 1711.920 ;
  LAYER metal4 ;
  RECT 1490.880 1710.800 1494.420 1711.920 ;
  LAYER metal3 ;
  RECT 1490.880 1710.800 1494.420 1711.920 ;
  LAYER metal2 ;
  RECT 1490.880 1710.800 1494.420 1711.920 ;
  LAYER metal1 ;
  RECT 1490.880 1710.800 1494.420 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1482.200 1710.800 1485.740 1711.920 ;
  LAYER metal4 ;
  RECT 1482.200 1710.800 1485.740 1711.920 ;
  LAYER metal3 ;
  RECT 1482.200 1710.800 1485.740 1711.920 ;
  LAYER metal2 ;
  RECT 1482.200 1710.800 1485.740 1711.920 ;
  LAYER metal1 ;
  RECT 1482.200 1710.800 1485.740 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1473.520 1710.800 1477.060 1711.920 ;
  LAYER metal4 ;
  RECT 1473.520 1710.800 1477.060 1711.920 ;
  LAYER metal3 ;
  RECT 1473.520 1710.800 1477.060 1711.920 ;
  LAYER metal2 ;
  RECT 1473.520 1710.800 1477.060 1711.920 ;
  LAYER metal1 ;
  RECT 1473.520 1710.800 1477.060 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1430.120 1710.800 1433.660 1711.920 ;
  LAYER metal4 ;
  RECT 1430.120 1710.800 1433.660 1711.920 ;
  LAYER metal3 ;
  RECT 1430.120 1710.800 1433.660 1711.920 ;
  LAYER metal2 ;
  RECT 1430.120 1710.800 1433.660 1711.920 ;
  LAYER metal1 ;
  RECT 1430.120 1710.800 1433.660 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1421.440 1710.800 1424.980 1711.920 ;
  LAYER metal4 ;
  RECT 1421.440 1710.800 1424.980 1711.920 ;
  LAYER metal3 ;
  RECT 1421.440 1710.800 1424.980 1711.920 ;
  LAYER metal2 ;
  RECT 1421.440 1710.800 1424.980 1711.920 ;
  LAYER metal1 ;
  RECT 1421.440 1710.800 1424.980 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1412.760 1710.800 1416.300 1711.920 ;
  LAYER metal4 ;
  RECT 1412.760 1710.800 1416.300 1711.920 ;
  LAYER metal3 ;
  RECT 1412.760 1710.800 1416.300 1711.920 ;
  LAYER metal2 ;
  RECT 1412.760 1710.800 1416.300 1711.920 ;
  LAYER metal1 ;
  RECT 1412.760 1710.800 1416.300 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1404.080 1710.800 1407.620 1711.920 ;
  LAYER metal4 ;
  RECT 1404.080 1710.800 1407.620 1711.920 ;
  LAYER metal3 ;
  RECT 1404.080 1710.800 1407.620 1711.920 ;
  LAYER metal2 ;
  RECT 1404.080 1710.800 1407.620 1711.920 ;
  LAYER metal1 ;
  RECT 1404.080 1710.800 1407.620 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1395.400 1710.800 1398.940 1711.920 ;
  LAYER metal4 ;
  RECT 1395.400 1710.800 1398.940 1711.920 ;
  LAYER metal3 ;
  RECT 1395.400 1710.800 1398.940 1711.920 ;
  LAYER metal2 ;
  RECT 1395.400 1710.800 1398.940 1711.920 ;
  LAYER metal1 ;
  RECT 1395.400 1710.800 1398.940 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1386.720 1710.800 1390.260 1711.920 ;
  LAYER metal4 ;
  RECT 1386.720 1710.800 1390.260 1711.920 ;
  LAYER metal3 ;
  RECT 1386.720 1710.800 1390.260 1711.920 ;
  LAYER metal2 ;
  RECT 1386.720 1710.800 1390.260 1711.920 ;
  LAYER metal1 ;
  RECT 1386.720 1710.800 1390.260 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1338.980 1710.800 1342.520 1711.920 ;
  LAYER metal4 ;
  RECT 1338.980 1710.800 1342.520 1711.920 ;
  LAYER metal3 ;
  RECT 1338.980 1710.800 1342.520 1711.920 ;
  LAYER metal2 ;
  RECT 1338.980 1710.800 1342.520 1711.920 ;
  LAYER metal1 ;
  RECT 1338.980 1710.800 1342.520 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1325.340 1710.800 1328.880 1711.920 ;
  LAYER metal4 ;
  RECT 1325.340 1710.800 1328.880 1711.920 ;
  LAYER metal3 ;
  RECT 1325.340 1710.800 1328.880 1711.920 ;
  LAYER metal2 ;
  RECT 1325.340 1710.800 1328.880 1711.920 ;
  LAYER metal1 ;
  RECT 1325.340 1710.800 1328.880 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1311.700 1710.800 1315.240 1711.920 ;
  LAYER metal4 ;
  RECT 1311.700 1710.800 1315.240 1711.920 ;
  LAYER metal3 ;
  RECT 1311.700 1710.800 1315.240 1711.920 ;
  LAYER metal2 ;
  RECT 1311.700 1710.800 1315.240 1711.920 ;
  LAYER metal1 ;
  RECT 1311.700 1710.800 1315.240 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1297.440 1710.800 1300.980 1711.920 ;
  LAYER metal4 ;
  RECT 1297.440 1710.800 1300.980 1711.920 ;
  LAYER metal3 ;
  RECT 1297.440 1710.800 1300.980 1711.920 ;
  LAYER metal2 ;
  RECT 1297.440 1710.800 1300.980 1711.920 ;
  LAYER metal1 ;
  RECT 1297.440 1710.800 1300.980 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1288.760 1710.800 1292.300 1711.920 ;
  LAYER metal4 ;
  RECT 1288.760 1710.800 1292.300 1711.920 ;
  LAYER metal3 ;
  RECT 1288.760 1710.800 1292.300 1711.920 ;
  LAYER metal2 ;
  RECT 1288.760 1710.800 1292.300 1711.920 ;
  LAYER metal1 ;
  RECT 1288.760 1710.800 1292.300 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1280.080 1710.800 1283.620 1711.920 ;
  LAYER metal4 ;
  RECT 1280.080 1710.800 1283.620 1711.920 ;
  LAYER metal3 ;
  RECT 1280.080 1710.800 1283.620 1711.920 ;
  LAYER metal2 ;
  RECT 1280.080 1710.800 1283.620 1711.920 ;
  LAYER metal1 ;
  RECT 1280.080 1710.800 1283.620 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1236.680 1710.800 1240.220 1711.920 ;
  LAYER metal4 ;
  RECT 1236.680 1710.800 1240.220 1711.920 ;
  LAYER metal3 ;
  RECT 1236.680 1710.800 1240.220 1711.920 ;
  LAYER metal2 ;
  RECT 1236.680 1710.800 1240.220 1711.920 ;
  LAYER metal1 ;
  RECT 1236.680 1710.800 1240.220 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1228.000 1710.800 1231.540 1711.920 ;
  LAYER metal4 ;
  RECT 1228.000 1710.800 1231.540 1711.920 ;
  LAYER metal3 ;
  RECT 1228.000 1710.800 1231.540 1711.920 ;
  LAYER metal2 ;
  RECT 1228.000 1710.800 1231.540 1711.920 ;
  LAYER metal1 ;
  RECT 1228.000 1710.800 1231.540 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1219.320 1710.800 1222.860 1711.920 ;
  LAYER metal4 ;
  RECT 1219.320 1710.800 1222.860 1711.920 ;
  LAYER metal3 ;
  RECT 1219.320 1710.800 1222.860 1711.920 ;
  LAYER metal2 ;
  RECT 1219.320 1710.800 1222.860 1711.920 ;
  LAYER metal1 ;
  RECT 1219.320 1710.800 1222.860 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1210.640 1710.800 1214.180 1711.920 ;
  LAYER metal4 ;
  RECT 1210.640 1710.800 1214.180 1711.920 ;
  LAYER metal3 ;
  RECT 1210.640 1710.800 1214.180 1711.920 ;
  LAYER metal2 ;
  RECT 1210.640 1710.800 1214.180 1711.920 ;
  LAYER metal1 ;
  RECT 1210.640 1710.800 1214.180 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1201.960 1710.800 1205.500 1711.920 ;
  LAYER metal4 ;
  RECT 1201.960 1710.800 1205.500 1711.920 ;
  LAYER metal3 ;
  RECT 1201.960 1710.800 1205.500 1711.920 ;
  LAYER metal2 ;
  RECT 1201.960 1710.800 1205.500 1711.920 ;
  LAYER metal1 ;
  RECT 1201.960 1710.800 1205.500 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1193.280 1710.800 1196.820 1711.920 ;
  LAYER metal4 ;
  RECT 1193.280 1710.800 1196.820 1711.920 ;
  LAYER metal3 ;
  RECT 1193.280 1710.800 1196.820 1711.920 ;
  LAYER metal2 ;
  RECT 1193.280 1710.800 1196.820 1711.920 ;
  LAYER metal1 ;
  RECT 1193.280 1710.800 1196.820 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1149.880 1710.800 1153.420 1711.920 ;
  LAYER metal4 ;
  RECT 1149.880 1710.800 1153.420 1711.920 ;
  LAYER metal3 ;
  RECT 1149.880 1710.800 1153.420 1711.920 ;
  LAYER metal2 ;
  RECT 1149.880 1710.800 1153.420 1711.920 ;
  LAYER metal1 ;
  RECT 1149.880 1710.800 1153.420 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1141.200 1710.800 1144.740 1711.920 ;
  LAYER metal4 ;
  RECT 1141.200 1710.800 1144.740 1711.920 ;
  LAYER metal3 ;
  RECT 1141.200 1710.800 1144.740 1711.920 ;
  LAYER metal2 ;
  RECT 1141.200 1710.800 1144.740 1711.920 ;
  LAYER metal1 ;
  RECT 1141.200 1710.800 1144.740 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1132.520 1710.800 1136.060 1711.920 ;
  LAYER metal4 ;
  RECT 1132.520 1710.800 1136.060 1711.920 ;
  LAYER metal3 ;
  RECT 1132.520 1710.800 1136.060 1711.920 ;
  LAYER metal2 ;
  RECT 1132.520 1710.800 1136.060 1711.920 ;
  LAYER metal1 ;
  RECT 1132.520 1710.800 1136.060 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1123.840 1710.800 1127.380 1711.920 ;
  LAYER metal4 ;
  RECT 1123.840 1710.800 1127.380 1711.920 ;
  LAYER metal3 ;
  RECT 1123.840 1710.800 1127.380 1711.920 ;
  LAYER metal2 ;
  RECT 1123.840 1710.800 1127.380 1711.920 ;
  LAYER metal1 ;
  RECT 1123.840 1710.800 1127.380 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1115.160 1710.800 1118.700 1711.920 ;
  LAYER metal4 ;
  RECT 1115.160 1710.800 1118.700 1711.920 ;
  LAYER metal3 ;
  RECT 1115.160 1710.800 1118.700 1711.920 ;
  LAYER metal2 ;
  RECT 1115.160 1710.800 1118.700 1711.920 ;
  LAYER metal1 ;
  RECT 1115.160 1710.800 1118.700 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1106.480 1710.800 1110.020 1711.920 ;
  LAYER metal4 ;
  RECT 1106.480 1710.800 1110.020 1711.920 ;
  LAYER metal3 ;
  RECT 1106.480 1710.800 1110.020 1711.920 ;
  LAYER metal2 ;
  RECT 1106.480 1710.800 1110.020 1711.920 ;
  LAYER metal1 ;
  RECT 1106.480 1710.800 1110.020 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1063.080 1710.800 1066.620 1711.920 ;
  LAYER metal4 ;
  RECT 1063.080 1710.800 1066.620 1711.920 ;
  LAYER metal3 ;
  RECT 1063.080 1710.800 1066.620 1711.920 ;
  LAYER metal2 ;
  RECT 1063.080 1710.800 1066.620 1711.920 ;
  LAYER metal1 ;
  RECT 1063.080 1710.800 1066.620 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1054.400 1710.800 1057.940 1711.920 ;
  LAYER metal4 ;
  RECT 1054.400 1710.800 1057.940 1711.920 ;
  LAYER metal3 ;
  RECT 1054.400 1710.800 1057.940 1711.920 ;
  LAYER metal2 ;
  RECT 1054.400 1710.800 1057.940 1711.920 ;
  LAYER metal1 ;
  RECT 1054.400 1710.800 1057.940 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1045.720 1710.800 1049.260 1711.920 ;
  LAYER metal4 ;
  RECT 1045.720 1710.800 1049.260 1711.920 ;
  LAYER metal3 ;
  RECT 1045.720 1710.800 1049.260 1711.920 ;
  LAYER metal2 ;
  RECT 1045.720 1710.800 1049.260 1711.920 ;
  LAYER metal1 ;
  RECT 1045.720 1710.800 1049.260 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1037.040 1710.800 1040.580 1711.920 ;
  LAYER metal4 ;
  RECT 1037.040 1710.800 1040.580 1711.920 ;
  LAYER metal3 ;
  RECT 1037.040 1710.800 1040.580 1711.920 ;
  LAYER metal2 ;
  RECT 1037.040 1710.800 1040.580 1711.920 ;
  LAYER metal1 ;
  RECT 1037.040 1710.800 1040.580 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1028.360 1710.800 1031.900 1711.920 ;
  LAYER metal4 ;
  RECT 1028.360 1710.800 1031.900 1711.920 ;
  LAYER metal3 ;
  RECT 1028.360 1710.800 1031.900 1711.920 ;
  LAYER metal2 ;
  RECT 1028.360 1710.800 1031.900 1711.920 ;
  LAYER metal1 ;
  RECT 1028.360 1710.800 1031.900 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1019.680 1710.800 1023.220 1711.920 ;
  LAYER metal4 ;
  RECT 1019.680 1710.800 1023.220 1711.920 ;
  LAYER metal3 ;
  RECT 1019.680 1710.800 1023.220 1711.920 ;
  LAYER metal2 ;
  RECT 1019.680 1710.800 1023.220 1711.920 ;
  LAYER metal1 ;
  RECT 1019.680 1710.800 1023.220 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 976.280 1710.800 979.820 1711.920 ;
  LAYER metal4 ;
  RECT 976.280 1710.800 979.820 1711.920 ;
  LAYER metal3 ;
  RECT 976.280 1710.800 979.820 1711.920 ;
  LAYER metal2 ;
  RECT 976.280 1710.800 979.820 1711.920 ;
  LAYER metal1 ;
  RECT 976.280 1710.800 979.820 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 967.600 1710.800 971.140 1711.920 ;
  LAYER metal4 ;
  RECT 967.600 1710.800 971.140 1711.920 ;
  LAYER metal3 ;
  RECT 967.600 1710.800 971.140 1711.920 ;
  LAYER metal2 ;
  RECT 967.600 1710.800 971.140 1711.920 ;
  LAYER metal1 ;
  RECT 967.600 1710.800 971.140 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 958.920 1710.800 962.460 1711.920 ;
  LAYER metal4 ;
  RECT 958.920 1710.800 962.460 1711.920 ;
  LAYER metal3 ;
  RECT 958.920 1710.800 962.460 1711.920 ;
  LAYER metal2 ;
  RECT 958.920 1710.800 962.460 1711.920 ;
  LAYER metal1 ;
  RECT 958.920 1710.800 962.460 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 950.240 1710.800 953.780 1711.920 ;
  LAYER metal4 ;
  RECT 950.240 1710.800 953.780 1711.920 ;
  LAYER metal3 ;
  RECT 950.240 1710.800 953.780 1711.920 ;
  LAYER metal2 ;
  RECT 950.240 1710.800 953.780 1711.920 ;
  LAYER metal1 ;
  RECT 950.240 1710.800 953.780 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 941.560 1710.800 945.100 1711.920 ;
  LAYER metal4 ;
  RECT 941.560 1710.800 945.100 1711.920 ;
  LAYER metal3 ;
  RECT 941.560 1710.800 945.100 1711.920 ;
  LAYER metal2 ;
  RECT 941.560 1710.800 945.100 1711.920 ;
  LAYER metal1 ;
  RECT 941.560 1710.800 945.100 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 932.880 1710.800 936.420 1711.920 ;
  LAYER metal4 ;
  RECT 932.880 1710.800 936.420 1711.920 ;
  LAYER metal3 ;
  RECT 932.880 1710.800 936.420 1711.920 ;
  LAYER metal2 ;
  RECT 932.880 1710.800 936.420 1711.920 ;
  LAYER metal1 ;
  RECT 932.880 1710.800 936.420 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 869.640 1710.800 873.180 1711.920 ;
  LAYER metal4 ;
  RECT 869.640 1710.800 873.180 1711.920 ;
  LAYER metal3 ;
  RECT 869.640 1710.800 873.180 1711.920 ;
  LAYER metal2 ;
  RECT 869.640 1710.800 873.180 1711.920 ;
  LAYER metal1 ;
  RECT 869.640 1710.800 873.180 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 860.960 1710.800 864.500 1711.920 ;
  LAYER metal4 ;
  RECT 860.960 1710.800 864.500 1711.920 ;
  LAYER metal3 ;
  RECT 860.960 1710.800 864.500 1711.920 ;
  LAYER metal2 ;
  RECT 860.960 1710.800 864.500 1711.920 ;
  LAYER metal1 ;
  RECT 860.960 1710.800 864.500 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 852.280 1710.800 855.820 1711.920 ;
  LAYER metal4 ;
  RECT 852.280 1710.800 855.820 1711.920 ;
  LAYER metal3 ;
  RECT 852.280 1710.800 855.820 1711.920 ;
  LAYER metal2 ;
  RECT 852.280 1710.800 855.820 1711.920 ;
  LAYER metal1 ;
  RECT 852.280 1710.800 855.820 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 843.600 1710.800 847.140 1711.920 ;
  LAYER metal4 ;
  RECT 843.600 1710.800 847.140 1711.920 ;
  LAYER metal3 ;
  RECT 843.600 1710.800 847.140 1711.920 ;
  LAYER metal2 ;
  RECT 843.600 1710.800 847.140 1711.920 ;
  LAYER metal1 ;
  RECT 843.600 1710.800 847.140 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 834.920 1710.800 838.460 1711.920 ;
  LAYER metal4 ;
  RECT 834.920 1710.800 838.460 1711.920 ;
  LAYER metal3 ;
  RECT 834.920 1710.800 838.460 1711.920 ;
  LAYER metal2 ;
  RECT 834.920 1710.800 838.460 1711.920 ;
  LAYER metal1 ;
  RECT 834.920 1710.800 838.460 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 826.240 1710.800 829.780 1711.920 ;
  LAYER metal4 ;
  RECT 826.240 1710.800 829.780 1711.920 ;
  LAYER metal3 ;
  RECT 826.240 1710.800 829.780 1711.920 ;
  LAYER metal2 ;
  RECT 826.240 1710.800 829.780 1711.920 ;
  LAYER metal1 ;
  RECT 826.240 1710.800 829.780 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 782.840 1710.800 786.380 1711.920 ;
  LAYER metal4 ;
  RECT 782.840 1710.800 786.380 1711.920 ;
  LAYER metal3 ;
  RECT 782.840 1710.800 786.380 1711.920 ;
  LAYER metal2 ;
  RECT 782.840 1710.800 786.380 1711.920 ;
  LAYER metal1 ;
  RECT 782.840 1710.800 786.380 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 774.160 1710.800 777.700 1711.920 ;
  LAYER metal4 ;
  RECT 774.160 1710.800 777.700 1711.920 ;
  LAYER metal3 ;
  RECT 774.160 1710.800 777.700 1711.920 ;
  LAYER metal2 ;
  RECT 774.160 1710.800 777.700 1711.920 ;
  LAYER metal1 ;
  RECT 774.160 1710.800 777.700 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 765.480 1710.800 769.020 1711.920 ;
  LAYER metal4 ;
  RECT 765.480 1710.800 769.020 1711.920 ;
  LAYER metal3 ;
  RECT 765.480 1710.800 769.020 1711.920 ;
  LAYER metal2 ;
  RECT 765.480 1710.800 769.020 1711.920 ;
  LAYER metal1 ;
  RECT 765.480 1710.800 769.020 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 756.800 1710.800 760.340 1711.920 ;
  LAYER metal4 ;
  RECT 756.800 1710.800 760.340 1711.920 ;
  LAYER metal3 ;
  RECT 756.800 1710.800 760.340 1711.920 ;
  LAYER metal2 ;
  RECT 756.800 1710.800 760.340 1711.920 ;
  LAYER metal1 ;
  RECT 756.800 1710.800 760.340 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 748.120 1710.800 751.660 1711.920 ;
  LAYER metal4 ;
  RECT 748.120 1710.800 751.660 1711.920 ;
  LAYER metal3 ;
  RECT 748.120 1710.800 751.660 1711.920 ;
  LAYER metal2 ;
  RECT 748.120 1710.800 751.660 1711.920 ;
  LAYER metal1 ;
  RECT 748.120 1710.800 751.660 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 739.440 1710.800 742.980 1711.920 ;
  LAYER metal4 ;
  RECT 739.440 1710.800 742.980 1711.920 ;
  LAYER metal3 ;
  RECT 739.440 1710.800 742.980 1711.920 ;
  LAYER metal2 ;
  RECT 739.440 1710.800 742.980 1711.920 ;
  LAYER metal1 ;
  RECT 739.440 1710.800 742.980 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 696.040 1710.800 699.580 1711.920 ;
  LAYER metal4 ;
  RECT 696.040 1710.800 699.580 1711.920 ;
  LAYER metal3 ;
  RECT 696.040 1710.800 699.580 1711.920 ;
  LAYER metal2 ;
  RECT 696.040 1710.800 699.580 1711.920 ;
  LAYER metal1 ;
  RECT 696.040 1710.800 699.580 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 687.360 1710.800 690.900 1711.920 ;
  LAYER metal4 ;
  RECT 687.360 1710.800 690.900 1711.920 ;
  LAYER metal3 ;
  RECT 687.360 1710.800 690.900 1711.920 ;
  LAYER metal2 ;
  RECT 687.360 1710.800 690.900 1711.920 ;
  LAYER metal1 ;
  RECT 687.360 1710.800 690.900 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 678.680 1710.800 682.220 1711.920 ;
  LAYER metal4 ;
  RECT 678.680 1710.800 682.220 1711.920 ;
  LAYER metal3 ;
  RECT 678.680 1710.800 682.220 1711.920 ;
  LAYER metal2 ;
  RECT 678.680 1710.800 682.220 1711.920 ;
  LAYER metal1 ;
  RECT 678.680 1710.800 682.220 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 670.000 1710.800 673.540 1711.920 ;
  LAYER metal4 ;
  RECT 670.000 1710.800 673.540 1711.920 ;
  LAYER metal3 ;
  RECT 670.000 1710.800 673.540 1711.920 ;
  LAYER metal2 ;
  RECT 670.000 1710.800 673.540 1711.920 ;
  LAYER metal1 ;
  RECT 670.000 1710.800 673.540 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 661.320 1710.800 664.860 1711.920 ;
  LAYER metal4 ;
  RECT 661.320 1710.800 664.860 1711.920 ;
  LAYER metal3 ;
  RECT 661.320 1710.800 664.860 1711.920 ;
  LAYER metal2 ;
  RECT 661.320 1710.800 664.860 1711.920 ;
  LAYER metal1 ;
  RECT 661.320 1710.800 664.860 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 652.640 1710.800 656.180 1711.920 ;
  LAYER metal4 ;
  RECT 652.640 1710.800 656.180 1711.920 ;
  LAYER metal3 ;
  RECT 652.640 1710.800 656.180 1711.920 ;
  LAYER metal2 ;
  RECT 652.640 1710.800 656.180 1711.920 ;
  LAYER metal1 ;
  RECT 652.640 1710.800 656.180 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 609.240 1710.800 612.780 1711.920 ;
  LAYER metal4 ;
  RECT 609.240 1710.800 612.780 1711.920 ;
  LAYER metal3 ;
  RECT 609.240 1710.800 612.780 1711.920 ;
  LAYER metal2 ;
  RECT 609.240 1710.800 612.780 1711.920 ;
  LAYER metal1 ;
  RECT 609.240 1710.800 612.780 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 600.560 1710.800 604.100 1711.920 ;
  LAYER metal4 ;
  RECT 600.560 1710.800 604.100 1711.920 ;
  LAYER metal3 ;
  RECT 600.560 1710.800 604.100 1711.920 ;
  LAYER metal2 ;
  RECT 600.560 1710.800 604.100 1711.920 ;
  LAYER metal1 ;
  RECT 600.560 1710.800 604.100 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 591.880 1710.800 595.420 1711.920 ;
  LAYER metal4 ;
  RECT 591.880 1710.800 595.420 1711.920 ;
  LAYER metal3 ;
  RECT 591.880 1710.800 595.420 1711.920 ;
  LAYER metal2 ;
  RECT 591.880 1710.800 595.420 1711.920 ;
  LAYER metal1 ;
  RECT 591.880 1710.800 595.420 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 583.200 1710.800 586.740 1711.920 ;
  LAYER metal4 ;
  RECT 583.200 1710.800 586.740 1711.920 ;
  LAYER metal3 ;
  RECT 583.200 1710.800 586.740 1711.920 ;
  LAYER metal2 ;
  RECT 583.200 1710.800 586.740 1711.920 ;
  LAYER metal1 ;
  RECT 583.200 1710.800 586.740 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 574.520 1710.800 578.060 1711.920 ;
  LAYER metal4 ;
  RECT 574.520 1710.800 578.060 1711.920 ;
  LAYER metal3 ;
  RECT 574.520 1710.800 578.060 1711.920 ;
  LAYER metal2 ;
  RECT 574.520 1710.800 578.060 1711.920 ;
  LAYER metal1 ;
  RECT 574.520 1710.800 578.060 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 565.840 1710.800 569.380 1711.920 ;
  LAYER metal4 ;
  RECT 565.840 1710.800 569.380 1711.920 ;
  LAYER metal3 ;
  RECT 565.840 1710.800 569.380 1711.920 ;
  LAYER metal2 ;
  RECT 565.840 1710.800 569.380 1711.920 ;
  LAYER metal1 ;
  RECT 565.840 1710.800 569.380 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 522.440 1710.800 525.980 1711.920 ;
  LAYER metal4 ;
  RECT 522.440 1710.800 525.980 1711.920 ;
  LAYER metal3 ;
  RECT 522.440 1710.800 525.980 1711.920 ;
  LAYER metal2 ;
  RECT 522.440 1710.800 525.980 1711.920 ;
  LAYER metal1 ;
  RECT 522.440 1710.800 525.980 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 513.760 1710.800 517.300 1711.920 ;
  LAYER metal4 ;
  RECT 513.760 1710.800 517.300 1711.920 ;
  LAYER metal3 ;
  RECT 513.760 1710.800 517.300 1711.920 ;
  LAYER metal2 ;
  RECT 513.760 1710.800 517.300 1711.920 ;
  LAYER metal1 ;
  RECT 513.760 1710.800 517.300 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 505.080 1710.800 508.620 1711.920 ;
  LAYER metal4 ;
  RECT 505.080 1710.800 508.620 1711.920 ;
  LAYER metal3 ;
  RECT 505.080 1710.800 508.620 1711.920 ;
  LAYER metal2 ;
  RECT 505.080 1710.800 508.620 1711.920 ;
  LAYER metal1 ;
  RECT 505.080 1710.800 508.620 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 496.400 1710.800 499.940 1711.920 ;
  LAYER metal4 ;
  RECT 496.400 1710.800 499.940 1711.920 ;
  LAYER metal3 ;
  RECT 496.400 1710.800 499.940 1711.920 ;
  LAYER metal2 ;
  RECT 496.400 1710.800 499.940 1711.920 ;
  LAYER metal1 ;
  RECT 496.400 1710.800 499.940 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 487.720 1710.800 491.260 1711.920 ;
  LAYER metal4 ;
  RECT 487.720 1710.800 491.260 1711.920 ;
  LAYER metal3 ;
  RECT 487.720 1710.800 491.260 1711.920 ;
  LAYER metal2 ;
  RECT 487.720 1710.800 491.260 1711.920 ;
  LAYER metal1 ;
  RECT 487.720 1710.800 491.260 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 474.080 1710.800 477.620 1711.920 ;
  LAYER metal4 ;
  RECT 474.080 1710.800 477.620 1711.920 ;
  LAYER metal3 ;
  RECT 474.080 1710.800 477.620 1711.920 ;
  LAYER metal2 ;
  RECT 474.080 1710.800 477.620 1711.920 ;
  LAYER metal1 ;
  RECT 474.080 1710.800 477.620 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 415.180 1710.800 418.720 1711.920 ;
  LAYER metal4 ;
  RECT 415.180 1710.800 418.720 1711.920 ;
  LAYER metal3 ;
  RECT 415.180 1710.800 418.720 1711.920 ;
  LAYER metal2 ;
  RECT 415.180 1710.800 418.720 1711.920 ;
  LAYER metal1 ;
  RECT 415.180 1710.800 418.720 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 406.500 1710.800 410.040 1711.920 ;
  LAYER metal4 ;
  RECT 406.500 1710.800 410.040 1711.920 ;
  LAYER metal3 ;
  RECT 406.500 1710.800 410.040 1711.920 ;
  LAYER metal2 ;
  RECT 406.500 1710.800 410.040 1711.920 ;
  LAYER metal1 ;
  RECT 406.500 1710.800 410.040 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 397.820 1710.800 401.360 1711.920 ;
  LAYER metal4 ;
  RECT 397.820 1710.800 401.360 1711.920 ;
  LAYER metal3 ;
  RECT 397.820 1710.800 401.360 1711.920 ;
  LAYER metal2 ;
  RECT 397.820 1710.800 401.360 1711.920 ;
  LAYER metal1 ;
  RECT 397.820 1710.800 401.360 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 389.140 1710.800 392.680 1711.920 ;
  LAYER metal4 ;
  RECT 389.140 1710.800 392.680 1711.920 ;
  LAYER metal3 ;
  RECT 389.140 1710.800 392.680 1711.920 ;
  LAYER metal2 ;
  RECT 389.140 1710.800 392.680 1711.920 ;
  LAYER metal1 ;
  RECT 389.140 1710.800 392.680 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 380.460 1710.800 384.000 1711.920 ;
  LAYER metal4 ;
  RECT 380.460 1710.800 384.000 1711.920 ;
  LAYER metal3 ;
  RECT 380.460 1710.800 384.000 1711.920 ;
  LAYER metal2 ;
  RECT 380.460 1710.800 384.000 1711.920 ;
  LAYER metal1 ;
  RECT 380.460 1710.800 384.000 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 371.780 1710.800 375.320 1711.920 ;
  LAYER metal4 ;
  RECT 371.780 1710.800 375.320 1711.920 ;
  LAYER metal3 ;
  RECT 371.780 1710.800 375.320 1711.920 ;
  LAYER metal2 ;
  RECT 371.780 1710.800 375.320 1711.920 ;
  LAYER metal1 ;
  RECT 371.780 1710.800 375.320 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 328.380 1710.800 331.920 1711.920 ;
  LAYER metal4 ;
  RECT 328.380 1710.800 331.920 1711.920 ;
  LAYER metal3 ;
  RECT 328.380 1710.800 331.920 1711.920 ;
  LAYER metal2 ;
  RECT 328.380 1710.800 331.920 1711.920 ;
  LAYER metal1 ;
  RECT 328.380 1710.800 331.920 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 319.700 1710.800 323.240 1711.920 ;
  LAYER metal4 ;
  RECT 319.700 1710.800 323.240 1711.920 ;
  LAYER metal3 ;
  RECT 319.700 1710.800 323.240 1711.920 ;
  LAYER metal2 ;
  RECT 319.700 1710.800 323.240 1711.920 ;
  LAYER metal1 ;
  RECT 319.700 1710.800 323.240 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 311.020 1710.800 314.560 1711.920 ;
  LAYER metal4 ;
  RECT 311.020 1710.800 314.560 1711.920 ;
  LAYER metal3 ;
  RECT 311.020 1710.800 314.560 1711.920 ;
  LAYER metal2 ;
  RECT 311.020 1710.800 314.560 1711.920 ;
  LAYER metal1 ;
  RECT 311.020 1710.800 314.560 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 302.340 1710.800 305.880 1711.920 ;
  LAYER metal4 ;
  RECT 302.340 1710.800 305.880 1711.920 ;
  LAYER metal3 ;
  RECT 302.340 1710.800 305.880 1711.920 ;
  LAYER metal2 ;
  RECT 302.340 1710.800 305.880 1711.920 ;
  LAYER metal1 ;
  RECT 302.340 1710.800 305.880 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 293.660 1710.800 297.200 1711.920 ;
  LAYER metal4 ;
  RECT 293.660 1710.800 297.200 1711.920 ;
  LAYER metal3 ;
  RECT 293.660 1710.800 297.200 1711.920 ;
  LAYER metal2 ;
  RECT 293.660 1710.800 297.200 1711.920 ;
  LAYER metal1 ;
  RECT 293.660 1710.800 297.200 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 284.980 1710.800 288.520 1711.920 ;
  LAYER metal4 ;
  RECT 284.980 1710.800 288.520 1711.920 ;
  LAYER metal3 ;
  RECT 284.980 1710.800 288.520 1711.920 ;
  LAYER metal2 ;
  RECT 284.980 1710.800 288.520 1711.920 ;
  LAYER metal1 ;
  RECT 284.980 1710.800 288.520 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 241.580 1710.800 245.120 1711.920 ;
  LAYER metal4 ;
  RECT 241.580 1710.800 245.120 1711.920 ;
  LAYER metal3 ;
  RECT 241.580 1710.800 245.120 1711.920 ;
  LAYER metal2 ;
  RECT 241.580 1710.800 245.120 1711.920 ;
  LAYER metal1 ;
  RECT 241.580 1710.800 245.120 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 232.900 1710.800 236.440 1711.920 ;
  LAYER metal4 ;
  RECT 232.900 1710.800 236.440 1711.920 ;
  LAYER metal3 ;
  RECT 232.900 1710.800 236.440 1711.920 ;
  LAYER metal2 ;
  RECT 232.900 1710.800 236.440 1711.920 ;
  LAYER metal1 ;
  RECT 232.900 1710.800 236.440 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 224.220 1710.800 227.760 1711.920 ;
  LAYER metal4 ;
  RECT 224.220 1710.800 227.760 1711.920 ;
  LAYER metal3 ;
  RECT 224.220 1710.800 227.760 1711.920 ;
  LAYER metal2 ;
  RECT 224.220 1710.800 227.760 1711.920 ;
  LAYER metal1 ;
  RECT 224.220 1710.800 227.760 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 215.540 1710.800 219.080 1711.920 ;
  LAYER metal4 ;
  RECT 215.540 1710.800 219.080 1711.920 ;
  LAYER metal3 ;
  RECT 215.540 1710.800 219.080 1711.920 ;
  LAYER metal2 ;
  RECT 215.540 1710.800 219.080 1711.920 ;
  LAYER metal1 ;
  RECT 215.540 1710.800 219.080 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 206.860 1710.800 210.400 1711.920 ;
  LAYER metal4 ;
  RECT 206.860 1710.800 210.400 1711.920 ;
  LAYER metal3 ;
  RECT 206.860 1710.800 210.400 1711.920 ;
  LAYER metal2 ;
  RECT 206.860 1710.800 210.400 1711.920 ;
  LAYER metal1 ;
  RECT 206.860 1710.800 210.400 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 198.180 1710.800 201.720 1711.920 ;
  LAYER metal4 ;
  RECT 198.180 1710.800 201.720 1711.920 ;
  LAYER metal3 ;
  RECT 198.180 1710.800 201.720 1711.920 ;
  LAYER metal2 ;
  RECT 198.180 1710.800 201.720 1711.920 ;
  LAYER metal1 ;
  RECT 198.180 1710.800 201.720 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 154.780 1710.800 158.320 1711.920 ;
  LAYER metal4 ;
  RECT 154.780 1710.800 158.320 1711.920 ;
  LAYER metal3 ;
  RECT 154.780 1710.800 158.320 1711.920 ;
  LAYER metal2 ;
  RECT 154.780 1710.800 158.320 1711.920 ;
  LAYER metal1 ;
  RECT 154.780 1710.800 158.320 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 146.100 1710.800 149.640 1711.920 ;
  LAYER metal4 ;
  RECT 146.100 1710.800 149.640 1711.920 ;
  LAYER metal3 ;
  RECT 146.100 1710.800 149.640 1711.920 ;
  LAYER metal2 ;
  RECT 146.100 1710.800 149.640 1711.920 ;
  LAYER metal1 ;
  RECT 146.100 1710.800 149.640 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 137.420 1710.800 140.960 1711.920 ;
  LAYER metal4 ;
  RECT 137.420 1710.800 140.960 1711.920 ;
  LAYER metal3 ;
  RECT 137.420 1710.800 140.960 1711.920 ;
  LAYER metal2 ;
  RECT 137.420 1710.800 140.960 1711.920 ;
  LAYER metal1 ;
  RECT 137.420 1710.800 140.960 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 128.740 1710.800 132.280 1711.920 ;
  LAYER metal4 ;
  RECT 128.740 1710.800 132.280 1711.920 ;
  LAYER metal3 ;
  RECT 128.740 1710.800 132.280 1711.920 ;
  LAYER metal2 ;
  RECT 128.740 1710.800 132.280 1711.920 ;
  LAYER metal1 ;
  RECT 128.740 1710.800 132.280 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 120.060 1710.800 123.600 1711.920 ;
  LAYER metal4 ;
  RECT 120.060 1710.800 123.600 1711.920 ;
  LAYER metal3 ;
  RECT 120.060 1710.800 123.600 1711.920 ;
  LAYER metal2 ;
  RECT 120.060 1710.800 123.600 1711.920 ;
  LAYER metal1 ;
  RECT 120.060 1710.800 123.600 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 111.380 1710.800 114.920 1711.920 ;
  LAYER metal4 ;
  RECT 111.380 1710.800 114.920 1711.920 ;
  LAYER metal3 ;
  RECT 111.380 1710.800 114.920 1711.920 ;
  LAYER metal2 ;
  RECT 111.380 1710.800 114.920 1711.920 ;
  LAYER metal1 ;
  RECT 111.380 1710.800 114.920 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 67.980 1710.800 71.520 1711.920 ;
  LAYER metal4 ;
  RECT 67.980 1710.800 71.520 1711.920 ;
  LAYER metal3 ;
  RECT 67.980 1710.800 71.520 1711.920 ;
  LAYER metal2 ;
  RECT 67.980 1710.800 71.520 1711.920 ;
  LAYER metal1 ;
  RECT 67.980 1710.800 71.520 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 59.300 1710.800 62.840 1711.920 ;
  LAYER metal4 ;
  RECT 59.300 1710.800 62.840 1711.920 ;
  LAYER metal3 ;
  RECT 59.300 1710.800 62.840 1711.920 ;
  LAYER metal2 ;
  RECT 59.300 1710.800 62.840 1711.920 ;
  LAYER metal1 ;
  RECT 59.300 1710.800 62.840 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 46.280 1710.800 49.820 1711.920 ;
  LAYER metal4 ;
  RECT 46.280 1710.800 49.820 1711.920 ;
  LAYER metal3 ;
  RECT 46.280 1710.800 49.820 1711.920 ;
  LAYER metal2 ;
  RECT 46.280 1710.800 49.820 1711.920 ;
  LAYER metal1 ;
  RECT 46.280 1710.800 49.820 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 32.640 1710.800 36.180 1711.920 ;
  LAYER metal4 ;
  RECT 32.640 1710.800 36.180 1711.920 ;
  LAYER metal3 ;
  RECT 32.640 1710.800 36.180 1711.920 ;
  LAYER metal2 ;
  RECT 32.640 1710.800 36.180 1711.920 ;
  LAYER metal1 ;
  RECT 32.640 1710.800 36.180 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 19.000 1710.800 22.540 1711.920 ;
  LAYER metal4 ;
  RECT 19.000 1710.800 22.540 1711.920 ;
  LAYER metal3 ;
  RECT 19.000 1710.800 22.540 1711.920 ;
  LAYER metal2 ;
  RECT 19.000 1710.800 22.540 1711.920 ;
  LAYER metal1 ;
  RECT 19.000 1710.800 22.540 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 7.220 1710.800 10.760 1711.920 ;
  LAYER metal4 ;
  RECT 7.220 1710.800 10.760 1711.920 ;
  LAYER metal3 ;
  RECT 7.220 1710.800 10.760 1711.920 ;
  LAYER metal2 ;
  RECT 7.220 1710.800 10.760 1711.920 ;
  LAYER metal1 ;
  RECT 7.220 1710.800 10.760 1711.920 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3587.720 0.000 3591.260 1.120 ;
  LAYER metal4 ;
  RECT 3587.720 0.000 3591.260 1.120 ;
  LAYER metal3 ;
  RECT 3587.720 0.000 3591.260 1.120 ;
  LAYER metal2 ;
  RECT 3587.720 0.000 3591.260 1.120 ;
  LAYER metal1 ;
  RECT 3587.720 0.000 3591.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3579.040 0.000 3582.580 1.120 ;
  LAYER metal4 ;
  RECT 3579.040 0.000 3582.580 1.120 ;
  LAYER metal3 ;
  RECT 3579.040 0.000 3582.580 1.120 ;
  LAYER metal2 ;
  RECT 3579.040 0.000 3582.580 1.120 ;
  LAYER metal1 ;
  RECT 3579.040 0.000 3582.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.360 0.000 3573.900 1.120 ;
  LAYER metal4 ;
  RECT 3570.360 0.000 3573.900 1.120 ;
  LAYER metal3 ;
  RECT 3570.360 0.000 3573.900 1.120 ;
  LAYER metal2 ;
  RECT 3570.360 0.000 3573.900 1.120 ;
  LAYER metal1 ;
  RECT 3570.360 0.000 3573.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3561.680 0.000 3565.220 1.120 ;
  LAYER metal4 ;
  RECT 3561.680 0.000 3565.220 1.120 ;
  LAYER metal3 ;
  RECT 3561.680 0.000 3565.220 1.120 ;
  LAYER metal2 ;
  RECT 3561.680 0.000 3565.220 1.120 ;
  LAYER metal1 ;
  RECT 3561.680 0.000 3565.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3553.000 0.000 3556.540 1.120 ;
  LAYER metal4 ;
  RECT 3553.000 0.000 3556.540 1.120 ;
  LAYER metal3 ;
  RECT 3553.000 0.000 3556.540 1.120 ;
  LAYER metal2 ;
  RECT 3553.000 0.000 3556.540 1.120 ;
  LAYER metal1 ;
  RECT 3553.000 0.000 3556.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3544.320 0.000 3547.860 1.120 ;
  LAYER metal4 ;
  RECT 3544.320 0.000 3547.860 1.120 ;
  LAYER metal3 ;
  RECT 3544.320 0.000 3547.860 1.120 ;
  LAYER metal2 ;
  RECT 3544.320 0.000 3547.860 1.120 ;
  LAYER metal1 ;
  RECT 3544.320 0.000 3547.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3500.920 0.000 3504.460 1.120 ;
  LAYER metal4 ;
  RECT 3500.920 0.000 3504.460 1.120 ;
  LAYER metal3 ;
  RECT 3500.920 0.000 3504.460 1.120 ;
  LAYER metal2 ;
  RECT 3500.920 0.000 3504.460 1.120 ;
  LAYER metal1 ;
  RECT 3500.920 0.000 3504.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3492.240 0.000 3495.780 1.120 ;
  LAYER metal4 ;
  RECT 3492.240 0.000 3495.780 1.120 ;
  LAYER metal3 ;
  RECT 3492.240 0.000 3495.780 1.120 ;
  LAYER metal2 ;
  RECT 3492.240 0.000 3495.780 1.120 ;
  LAYER metal1 ;
  RECT 3492.240 0.000 3495.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3483.560 0.000 3487.100 1.120 ;
  LAYER metal4 ;
  RECT 3483.560 0.000 3487.100 1.120 ;
  LAYER metal3 ;
  RECT 3483.560 0.000 3487.100 1.120 ;
  LAYER metal2 ;
  RECT 3483.560 0.000 3487.100 1.120 ;
  LAYER metal1 ;
  RECT 3483.560 0.000 3487.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3474.880 0.000 3478.420 1.120 ;
  LAYER metal4 ;
  RECT 3474.880 0.000 3478.420 1.120 ;
  LAYER metal3 ;
  RECT 3474.880 0.000 3478.420 1.120 ;
  LAYER metal2 ;
  RECT 3474.880 0.000 3478.420 1.120 ;
  LAYER metal1 ;
  RECT 3474.880 0.000 3478.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3466.200 0.000 3469.740 1.120 ;
  LAYER metal4 ;
  RECT 3466.200 0.000 3469.740 1.120 ;
  LAYER metal3 ;
  RECT 3466.200 0.000 3469.740 1.120 ;
  LAYER metal2 ;
  RECT 3466.200 0.000 3469.740 1.120 ;
  LAYER metal1 ;
  RECT 3466.200 0.000 3469.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3457.520 0.000 3461.060 1.120 ;
  LAYER metal4 ;
  RECT 3457.520 0.000 3461.060 1.120 ;
  LAYER metal3 ;
  RECT 3457.520 0.000 3461.060 1.120 ;
  LAYER metal2 ;
  RECT 3457.520 0.000 3461.060 1.120 ;
  LAYER metal1 ;
  RECT 3457.520 0.000 3461.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3414.120 0.000 3417.660 1.120 ;
  LAYER metal4 ;
  RECT 3414.120 0.000 3417.660 1.120 ;
  LAYER metal3 ;
  RECT 3414.120 0.000 3417.660 1.120 ;
  LAYER metal2 ;
  RECT 3414.120 0.000 3417.660 1.120 ;
  LAYER metal1 ;
  RECT 3414.120 0.000 3417.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3405.440 0.000 3408.980 1.120 ;
  LAYER metal4 ;
  RECT 3405.440 0.000 3408.980 1.120 ;
  LAYER metal3 ;
  RECT 3405.440 0.000 3408.980 1.120 ;
  LAYER metal2 ;
  RECT 3405.440 0.000 3408.980 1.120 ;
  LAYER metal1 ;
  RECT 3405.440 0.000 3408.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3396.760 0.000 3400.300 1.120 ;
  LAYER metal4 ;
  RECT 3396.760 0.000 3400.300 1.120 ;
  LAYER metal3 ;
  RECT 3396.760 0.000 3400.300 1.120 ;
  LAYER metal2 ;
  RECT 3396.760 0.000 3400.300 1.120 ;
  LAYER metal1 ;
  RECT 3396.760 0.000 3400.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3388.080 0.000 3391.620 1.120 ;
  LAYER metal4 ;
  RECT 3388.080 0.000 3391.620 1.120 ;
  LAYER metal3 ;
  RECT 3388.080 0.000 3391.620 1.120 ;
  LAYER metal2 ;
  RECT 3388.080 0.000 3391.620 1.120 ;
  LAYER metal1 ;
  RECT 3388.080 0.000 3391.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3379.400 0.000 3382.940 1.120 ;
  LAYER metal4 ;
  RECT 3379.400 0.000 3382.940 1.120 ;
  LAYER metal3 ;
  RECT 3379.400 0.000 3382.940 1.120 ;
  LAYER metal2 ;
  RECT 3379.400 0.000 3382.940 1.120 ;
  LAYER metal1 ;
  RECT 3379.400 0.000 3382.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3370.720 0.000 3374.260 1.120 ;
  LAYER metal4 ;
  RECT 3370.720 0.000 3374.260 1.120 ;
  LAYER metal3 ;
  RECT 3370.720 0.000 3374.260 1.120 ;
  LAYER metal2 ;
  RECT 3370.720 0.000 3374.260 1.120 ;
  LAYER metal1 ;
  RECT 3370.720 0.000 3374.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3327.320 0.000 3330.860 1.120 ;
  LAYER metal4 ;
  RECT 3327.320 0.000 3330.860 1.120 ;
  LAYER metal3 ;
  RECT 3327.320 0.000 3330.860 1.120 ;
  LAYER metal2 ;
  RECT 3327.320 0.000 3330.860 1.120 ;
  LAYER metal1 ;
  RECT 3327.320 0.000 3330.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3318.640 0.000 3322.180 1.120 ;
  LAYER metal4 ;
  RECT 3318.640 0.000 3322.180 1.120 ;
  LAYER metal3 ;
  RECT 3318.640 0.000 3322.180 1.120 ;
  LAYER metal2 ;
  RECT 3318.640 0.000 3322.180 1.120 ;
  LAYER metal1 ;
  RECT 3318.640 0.000 3322.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3309.960 0.000 3313.500 1.120 ;
  LAYER metal4 ;
  RECT 3309.960 0.000 3313.500 1.120 ;
  LAYER metal3 ;
  RECT 3309.960 0.000 3313.500 1.120 ;
  LAYER metal2 ;
  RECT 3309.960 0.000 3313.500 1.120 ;
  LAYER metal1 ;
  RECT 3309.960 0.000 3313.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3301.280 0.000 3304.820 1.120 ;
  LAYER metal4 ;
  RECT 3301.280 0.000 3304.820 1.120 ;
  LAYER metal3 ;
  RECT 3301.280 0.000 3304.820 1.120 ;
  LAYER metal2 ;
  RECT 3301.280 0.000 3304.820 1.120 ;
  LAYER metal1 ;
  RECT 3301.280 0.000 3304.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3292.600 0.000 3296.140 1.120 ;
  LAYER metal4 ;
  RECT 3292.600 0.000 3296.140 1.120 ;
  LAYER metal3 ;
  RECT 3292.600 0.000 3296.140 1.120 ;
  LAYER metal2 ;
  RECT 3292.600 0.000 3296.140 1.120 ;
  LAYER metal1 ;
  RECT 3292.600 0.000 3296.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3283.920 0.000 3287.460 1.120 ;
  LAYER metal4 ;
  RECT 3283.920 0.000 3287.460 1.120 ;
  LAYER metal3 ;
  RECT 3283.920 0.000 3287.460 1.120 ;
  LAYER metal2 ;
  RECT 3283.920 0.000 3287.460 1.120 ;
  LAYER metal1 ;
  RECT 3283.920 0.000 3287.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3240.520 0.000 3244.060 1.120 ;
  LAYER metal4 ;
  RECT 3240.520 0.000 3244.060 1.120 ;
  LAYER metal3 ;
  RECT 3240.520 0.000 3244.060 1.120 ;
  LAYER metal2 ;
  RECT 3240.520 0.000 3244.060 1.120 ;
  LAYER metal1 ;
  RECT 3240.520 0.000 3244.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3231.840 0.000 3235.380 1.120 ;
  LAYER metal4 ;
  RECT 3231.840 0.000 3235.380 1.120 ;
  LAYER metal3 ;
  RECT 3231.840 0.000 3235.380 1.120 ;
  LAYER metal2 ;
  RECT 3231.840 0.000 3235.380 1.120 ;
  LAYER metal1 ;
  RECT 3231.840 0.000 3235.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3223.160 0.000 3226.700 1.120 ;
  LAYER metal4 ;
  RECT 3223.160 0.000 3226.700 1.120 ;
  LAYER metal3 ;
  RECT 3223.160 0.000 3226.700 1.120 ;
  LAYER metal2 ;
  RECT 3223.160 0.000 3226.700 1.120 ;
  LAYER metal1 ;
  RECT 3223.160 0.000 3226.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3214.480 0.000 3218.020 1.120 ;
  LAYER metal4 ;
  RECT 3214.480 0.000 3218.020 1.120 ;
  LAYER metal3 ;
  RECT 3214.480 0.000 3218.020 1.120 ;
  LAYER metal2 ;
  RECT 3214.480 0.000 3218.020 1.120 ;
  LAYER metal1 ;
  RECT 3214.480 0.000 3218.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3201.460 0.000 3205.000 1.120 ;
  LAYER metal4 ;
  RECT 3201.460 0.000 3205.000 1.120 ;
  LAYER metal3 ;
  RECT 3201.460 0.000 3205.000 1.120 ;
  LAYER metal2 ;
  RECT 3201.460 0.000 3205.000 1.120 ;
  LAYER metal1 ;
  RECT 3201.460 0.000 3205.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3187.820 0.000 3191.360 1.120 ;
  LAYER metal4 ;
  RECT 3187.820 0.000 3191.360 1.120 ;
  LAYER metal3 ;
  RECT 3187.820 0.000 3191.360 1.120 ;
  LAYER metal2 ;
  RECT 3187.820 0.000 3191.360 1.120 ;
  LAYER metal1 ;
  RECT 3187.820 0.000 3191.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3133.880 0.000 3137.420 1.120 ;
  LAYER metal4 ;
  RECT 3133.880 0.000 3137.420 1.120 ;
  LAYER metal3 ;
  RECT 3133.880 0.000 3137.420 1.120 ;
  LAYER metal2 ;
  RECT 3133.880 0.000 3137.420 1.120 ;
  LAYER metal1 ;
  RECT 3133.880 0.000 3137.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3125.200 0.000 3128.740 1.120 ;
  LAYER metal4 ;
  RECT 3125.200 0.000 3128.740 1.120 ;
  LAYER metal3 ;
  RECT 3125.200 0.000 3128.740 1.120 ;
  LAYER metal2 ;
  RECT 3125.200 0.000 3128.740 1.120 ;
  LAYER metal1 ;
  RECT 3125.200 0.000 3128.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3116.520 0.000 3120.060 1.120 ;
  LAYER metal4 ;
  RECT 3116.520 0.000 3120.060 1.120 ;
  LAYER metal3 ;
  RECT 3116.520 0.000 3120.060 1.120 ;
  LAYER metal2 ;
  RECT 3116.520 0.000 3120.060 1.120 ;
  LAYER metal1 ;
  RECT 3116.520 0.000 3120.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3107.840 0.000 3111.380 1.120 ;
  LAYER metal4 ;
  RECT 3107.840 0.000 3111.380 1.120 ;
  LAYER metal3 ;
  RECT 3107.840 0.000 3111.380 1.120 ;
  LAYER metal2 ;
  RECT 3107.840 0.000 3111.380 1.120 ;
  LAYER metal1 ;
  RECT 3107.840 0.000 3111.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3099.160 0.000 3102.700 1.120 ;
  LAYER metal4 ;
  RECT 3099.160 0.000 3102.700 1.120 ;
  LAYER metal3 ;
  RECT 3099.160 0.000 3102.700 1.120 ;
  LAYER metal2 ;
  RECT 3099.160 0.000 3102.700 1.120 ;
  LAYER metal1 ;
  RECT 3099.160 0.000 3102.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3090.480 0.000 3094.020 1.120 ;
  LAYER metal4 ;
  RECT 3090.480 0.000 3094.020 1.120 ;
  LAYER metal3 ;
  RECT 3090.480 0.000 3094.020 1.120 ;
  LAYER metal2 ;
  RECT 3090.480 0.000 3094.020 1.120 ;
  LAYER metal1 ;
  RECT 3090.480 0.000 3094.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3047.080 0.000 3050.620 1.120 ;
  LAYER metal4 ;
  RECT 3047.080 0.000 3050.620 1.120 ;
  LAYER metal3 ;
  RECT 3047.080 0.000 3050.620 1.120 ;
  LAYER metal2 ;
  RECT 3047.080 0.000 3050.620 1.120 ;
  LAYER metal1 ;
  RECT 3047.080 0.000 3050.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3038.400 0.000 3041.940 1.120 ;
  LAYER metal4 ;
  RECT 3038.400 0.000 3041.940 1.120 ;
  LAYER metal3 ;
  RECT 3038.400 0.000 3041.940 1.120 ;
  LAYER metal2 ;
  RECT 3038.400 0.000 3041.940 1.120 ;
  LAYER metal1 ;
  RECT 3038.400 0.000 3041.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3029.720 0.000 3033.260 1.120 ;
  LAYER metal4 ;
  RECT 3029.720 0.000 3033.260 1.120 ;
  LAYER metal3 ;
  RECT 3029.720 0.000 3033.260 1.120 ;
  LAYER metal2 ;
  RECT 3029.720 0.000 3033.260 1.120 ;
  LAYER metal1 ;
  RECT 3029.720 0.000 3033.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3021.040 0.000 3024.580 1.120 ;
  LAYER metal4 ;
  RECT 3021.040 0.000 3024.580 1.120 ;
  LAYER metal3 ;
  RECT 3021.040 0.000 3024.580 1.120 ;
  LAYER metal2 ;
  RECT 3021.040 0.000 3024.580 1.120 ;
  LAYER metal1 ;
  RECT 3021.040 0.000 3024.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3012.360 0.000 3015.900 1.120 ;
  LAYER metal4 ;
  RECT 3012.360 0.000 3015.900 1.120 ;
  LAYER metal3 ;
  RECT 3012.360 0.000 3015.900 1.120 ;
  LAYER metal2 ;
  RECT 3012.360 0.000 3015.900 1.120 ;
  LAYER metal1 ;
  RECT 3012.360 0.000 3015.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3003.680 0.000 3007.220 1.120 ;
  LAYER metal4 ;
  RECT 3003.680 0.000 3007.220 1.120 ;
  LAYER metal3 ;
  RECT 3003.680 0.000 3007.220 1.120 ;
  LAYER metal2 ;
  RECT 3003.680 0.000 3007.220 1.120 ;
  LAYER metal1 ;
  RECT 3003.680 0.000 3007.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2960.280 0.000 2963.820 1.120 ;
  LAYER metal4 ;
  RECT 2960.280 0.000 2963.820 1.120 ;
  LAYER metal3 ;
  RECT 2960.280 0.000 2963.820 1.120 ;
  LAYER metal2 ;
  RECT 2960.280 0.000 2963.820 1.120 ;
  LAYER metal1 ;
  RECT 2960.280 0.000 2963.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2951.600 0.000 2955.140 1.120 ;
  LAYER metal4 ;
  RECT 2951.600 0.000 2955.140 1.120 ;
  LAYER metal3 ;
  RECT 2951.600 0.000 2955.140 1.120 ;
  LAYER metal2 ;
  RECT 2951.600 0.000 2955.140 1.120 ;
  LAYER metal1 ;
  RECT 2951.600 0.000 2955.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2942.920 0.000 2946.460 1.120 ;
  LAYER metal4 ;
  RECT 2942.920 0.000 2946.460 1.120 ;
  LAYER metal3 ;
  RECT 2942.920 0.000 2946.460 1.120 ;
  LAYER metal2 ;
  RECT 2942.920 0.000 2946.460 1.120 ;
  LAYER metal1 ;
  RECT 2942.920 0.000 2946.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2934.240 0.000 2937.780 1.120 ;
  LAYER metal4 ;
  RECT 2934.240 0.000 2937.780 1.120 ;
  LAYER metal3 ;
  RECT 2934.240 0.000 2937.780 1.120 ;
  LAYER metal2 ;
  RECT 2934.240 0.000 2937.780 1.120 ;
  LAYER metal1 ;
  RECT 2934.240 0.000 2937.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2925.560 0.000 2929.100 1.120 ;
  LAYER metal4 ;
  RECT 2925.560 0.000 2929.100 1.120 ;
  LAYER metal3 ;
  RECT 2925.560 0.000 2929.100 1.120 ;
  LAYER metal2 ;
  RECT 2925.560 0.000 2929.100 1.120 ;
  LAYER metal1 ;
  RECT 2925.560 0.000 2929.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2916.880 0.000 2920.420 1.120 ;
  LAYER metal4 ;
  RECT 2916.880 0.000 2920.420 1.120 ;
  LAYER metal3 ;
  RECT 2916.880 0.000 2920.420 1.120 ;
  LAYER metal2 ;
  RECT 2916.880 0.000 2920.420 1.120 ;
  LAYER metal1 ;
  RECT 2916.880 0.000 2920.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2873.480 0.000 2877.020 1.120 ;
  LAYER metal4 ;
  RECT 2873.480 0.000 2877.020 1.120 ;
  LAYER metal3 ;
  RECT 2873.480 0.000 2877.020 1.120 ;
  LAYER metal2 ;
  RECT 2873.480 0.000 2877.020 1.120 ;
  LAYER metal1 ;
  RECT 2873.480 0.000 2877.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2864.800 0.000 2868.340 1.120 ;
  LAYER metal4 ;
  RECT 2864.800 0.000 2868.340 1.120 ;
  LAYER metal3 ;
  RECT 2864.800 0.000 2868.340 1.120 ;
  LAYER metal2 ;
  RECT 2864.800 0.000 2868.340 1.120 ;
  LAYER metal1 ;
  RECT 2864.800 0.000 2868.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2856.120 0.000 2859.660 1.120 ;
  LAYER metal4 ;
  RECT 2856.120 0.000 2859.660 1.120 ;
  LAYER metal3 ;
  RECT 2856.120 0.000 2859.660 1.120 ;
  LAYER metal2 ;
  RECT 2856.120 0.000 2859.660 1.120 ;
  LAYER metal1 ;
  RECT 2856.120 0.000 2859.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2847.440 0.000 2850.980 1.120 ;
  LAYER metal4 ;
  RECT 2847.440 0.000 2850.980 1.120 ;
  LAYER metal3 ;
  RECT 2847.440 0.000 2850.980 1.120 ;
  LAYER metal2 ;
  RECT 2847.440 0.000 2850.980 1.120 ;
  LAYER metal1 ;
  RECT 2847.440 0.000 2850.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2838.760 0.000 2842.300 1.120 ;
  LAYER metal4 ;
  RECT 2838.760 0.000 2842.300 1.120 ;
  LAYER metal3 ;
  RECT 2838.760 0.000 2842.300 1.120 ;
  LAYER metal2 ;
  RECT 2838.760 0.000 2842.300 1.120 ;
  LAYER metal1 ;
  RECT 2838.760 0.000 2842.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2830.080 0.000 2833.620 1.120 ;
  LAYER metal4 ;
  RECT 2830.080 0.000 2833.620 1.120 ;
  LAYER metal3 ;
  RECT 2830.080 0.000 2833.620 1.120 ;
  LAYER metal2 ;
  RECT 2830.080 0.000 2833.620 1.120 ;
  LAYER metal1 ;
  RECT 2830.080 0.000 2833.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2786.680 0.000 2790.220 1.120 ;
  LAYER metal4 ;
  RECT 2786.680 0.000 2790.220 1.120 ;
  LAYER metal3 ;
  RECT 2786.680 0.000 2790.220 1.120 ;
  LAYER metal2 ;
  RECT 2786.680 0.000 2790.220 1.120 ;
  LAYER metal1 ;
  RECT 2786.680 0.000 2790.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2773.660 0.000 2777.200 1.120 ;
  LAYER metal4 ;
  RECT 2773.660 0.000 2777.200 1.120 ;
  LAYER metal3 ;
  RECT 2773.660 0.000 2777.200 1.120 ;
  LAYER metal2 ;
  RECT 2773.660 0.000 2777.200 1.120 ;
  LAYER metal1 ;
  RECT 2773.660 0.000 2777.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2760.020 0.000 2763.560 1.120 ;
  LAYER metal4 ;
  RECT 2760.020 0.000 2763.560 1.120 ;
  LAYER metal3 ;
  RECT 2760.020 0.000 2763.560 1.120 ;
  LAYER metal2 ;
  RECT 2760.020 0.000 2763.560 1.120 ;
  LAYER metal1 ;
  RECT 2760.020 0.000 2763.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2746.380 0.000 2749.920 1.120 ;
  LAYER metal4 ;
  RECT 2746.380 0.000 2749.920 1.120 ;
  LAYER metal3 ;
  RECT 2746.380 0.000 2749.920 1.120 ;
  LAYER metal2 ;
  RECT 2746.380 0.000 2749.920 1.120 ;
  LAYER metal1 ;
  RECT 2746.380 0.000 2749.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2732.120 0.000 2735.660 1.120 ;
  LAYER metal4 ;
  RECT 2732.120 0.000 2735.660 1.120 ;
  LAYER metal3 ;
  RECT 2732.120 0.000 2735.660 1.120 ;
  LAYER metal2 ;
  RECT 2732.120 0.000 2735.660 1.120 ;
  LAYER metal1 ;
  RECT 2732.120 0.000 2735.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2723.440 0.000 2726.980 1.120 ;
  LAYER metal4 ;
  RECT 2723.440 0.000 2726.980 1.120 ;
  LAYER metal3 ;
  RECT 2723.440 0.000 2726.980 1.120 ;
  LAYER metal2 ;
  RECT 2723.440 0.000 2726.980 1.120 ;
  LAYER metal1 ;
  RECT 2723.440 0.000 2726.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2680.040 0.000 2683.580 1.120 ;
  LAYER metal4 ;
  RECT 2680.040 0.000 2683.580 1.120 ;
  LAYER metal3 ;
  RECT 2680.040 0.000 2683.580 1.120 ;
  LAYER metal2 ;
  RECT 2680.040 0.000 2683.580 1.120 ;
  LAYER metal1 ;
  RECT 2680.040 0.000 2683.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2671.360 0.000 2674.900 1.120 ;
  LAYER metal4 ;
  RECT 2671.360 0.000 2674.900 1.120 ;
  LAYER metal3 ;
  RECT 2671.360 0.000 2674.900 1.120 ;
  LAYER metal2 ;
  RECT 2671.360 0.000 2674.900 1.120 ;
  LAYER metal1 ;
  RECT 2671.360 0.000 2674.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2662.680 0.000 2666.220 1.120 ;
  LAYER metal4 ;
  RECT 2662.680 0.000 2666.220 1.120 ;
  LAYER metal3 ;
  RECT 2662.680 0.000 2666.220 1.120 ;
  LAYER metal2 ;
  RECT 2662.680 0.000 2666.220 1.120 ;
  LAYER metal1 ;
  RECT 2662.680 0.000 2666.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2654.000 0.000 2657.540 1.120 ;
  LAYER metal4 ;
  RECT 2654.000 0.000 2657.540 1.120 ;
  LAYER metal3 ;
  RECT 2654.000 0.000 2657.540 1.120 ;
  LAYER metal2 ;
  RECT 2654.000 0.000 2657.540 1.120 ;
  LAYER metal1 ;
  RECT 2654.000 0.000 2657.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2645.320 0.000 2648.860 1.120 ;
  LAYER metal4 ;
  RECT 2645.320 0.000 2648.860 1.120 ;
  LAYER metal3 ;
  RECT 2645.320 0.000 2648.860 1.120 ;
  LAYER metal2 ;
  RECT 2645.320 0.000 2648.860 1.120 ;
  LAYER metal1 ;
  RECT 2645.320 0.000 2648.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2636.640 0.000 2640.180 1.120 ;
  LAYER metal4 ;
  RECT 2636.640 0.000 2640.180 1.120 ;
  LAYER metal3 ;
  RECT 2636.640 0.000 2640.180 1.120 ;
  LAYER metal2 ;
  RECT 2636.640 0.000 2640.180 1.120 ;
  LAYER metal1 ;
  RECT 2636.640 0.000 2640.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2593.240 0.000 2596.780 1.120 ;
  LAYER metal4 ;
  RECT 2593.240 0.000 2596.780 1.120 ;
  LAYER metal3 ;
  RECT 2593.240 0.000 2596.780 1.120 ;
  LAYER metal2 ;
  RECT 2593.240 0.000 2596.780 1.120 ;
  LAYER metal1 ;
  RECT 2593.240 0.000 2596.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2584.560 0.000 2588.100 1.120 ;
  LAYER metal4 ;
  RECT 2584.560 0.000 2588.100 1.120 ;
  LAYER metal3 ;
  RECT 2584.560 0.000 2588.100 1.120 ;
  LAYER metal2 ;
  RECT 2584.560 0.000 2588.100 1.120 ;
  LAYER metal1 ;
  RECT 2584.560 0.000 2588.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2575.880 0.000 2579.420 1.120 ;
  LAYER metal4 ;
  RECT 2575.880 0.000 2579.420 1.120 ;
  LAYER metal3 ;
  RECT 2575.880 0.000 2579.420 1.120 ;
  LAYER metal2 ;
  RECT 2575.880 0.000 2579.420 1.120 ;
  LAYER metal1 ;
  RECT 2575.880 0.000 2579.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2567.200 0.000 2570.740 1.120 ;
  LAYER metal4 ;
  RECT 2567.200 0.000 2570.740 1.120 ;
  LAYER metal3 ;
  RECT 2567.200 0.000 2570.740 1.120 ;
  LAYER metal2 ;
  RECT 2567.200 0.000 2570.740 1.120 ;
  LAYER metal1 ;
  RECT 2567.200 0.000 2570.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2558.520 0.000 2562.060 1.120 ;
  LAYER metal4 ;
  RECT 2558.520 0.000 2562.060 1.120 ;
  LAYER metal3 ;
  RECT 2558.520 0.000 2562.060 1.120 ;
  LAYER metal2 ;
  RECT 2558.520 0.000 2562.060 1.120 ;
  LAYER metal1 ;
  RECT 2558.520 0.000 2562.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2549.840 0.000 2553.380 1.120 ;
  LAYER metal4 ;
  RECT 2549.840 0.000 2553.380 1.120 ;
  LAYER metal3 ;
  RECT 2549.840 0.000 2553.380 1.120 ;
  LAYER metal2 ;
  RECT 2549.840 0.000 2553.380 1.120 ;
  LAYER metal1 ;
  RECT 2549.840 0.000 2553.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2506.440 0.000 2509.980 1.120 ;
  LAYER metal4 ;
  RECT 2506.440 0.000 2509.980 1.120 ;
  LAYER metal3 ;
  RECT 2506.440 0.000 2509.980 1.120 ;
  LAYER metal2 ;
  RECT 2506.440 0.000 2509.980 1.120 ;
  LAYER metal1 ;
  RECT 2506.440 0.000 2509.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2497.760 0.000 2501.300 1.120 ;
  LAYER metal4 ;
  RECT 2497.760 0.000 2501.300 1.120 ;
  LAYER metal3 ;
  RECT 2497.760 0.000 2501.300 1.120 ;
  LAYER metal2 ;
  RECT 2497.760 0.000 2501.300 1.120 ;
  LAYER metal1 ;
  RECT 2497.760 0.000 2501.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2489.080 0.000 2492.620 1.120 ;
  LAYER metal4 ;
  RECT 2489.080 0.000 2492.620 1.120 ;
  LAYER metal3 ;
  RECT 2489.080 0.000 2492.620 1.120 ;
  LAYER metal2 ;
  RECT 2489.080 0.000 2492.620 1.120 ;
  LAYER metal1 ;
  RECT 2489.080 0.000 2492.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2480.400 0.000 2483.940 1.120 ;
  LAYER metal4 ;
  RECT 2480.400 0.000 2483.940 1.120 ;
  LAYER metal3 ;
  RECT 2480.400 0.000 2483.940 1.120 ;
  LAYER metal2 ;
  RECT 2480.400 0.000 2483.940 1.120 ;
  LAYER metal1 ;
  RECT 2480.400 0.000 2483.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2471.720 0.000 2475.260 1.120 ;
  LAYER metal4 ;
  RECT 2471.720 0.000 2475.260 1.120 ;
  LAYER metal3 ;
  RECT 2471.720 0.000 2475.260 1.120 ;
  LAYER metal2 ;
  RECT 2471.720 0.000 2475.260 1.120 ;
  LAYER metal1 ;
  RECT 2471.720 0.000 2475.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2463.040 0.000 2466.580 1.120 ;
  LAYER metal4 ;
  RECT 2463.040 0.000 2466.580 1.120 ;
  LAYER metal3 ;
  RECT 2463.040 0.000 2466.580 1.120 ;
  LAYER metal2 ;
  RECT 2463.040 0.000 2466.580 1.120 ;
  LAYER metal1 ;
  RECT 2463.040 0.000 2466.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2419.640 0.000 2423.180 1.120 ;
  LAYER metal4 ;
  RECT 2419.640 0.000 2423.180 1.120 ;
  LAYER metal3 ;
  RECT 2419.640 0.000 2423.180 1.120 ;
  LAYER metal2 ;
  RECT 2419.640 0.000 2423.180 1.120 ;
  LAYER metal1 ;
  RECT 2419.640 0.000 2423.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2410.960 0.000 2414.500 1.120 ;
  LAYER metal4 ;
  RECT 2410.960 0.000 2414.500 1.120 ;
  LAYER metal3 ;
  RECT 2410.960 0.000 2414.500 1.120 ;
  LAYER metal2 ;
  RECT 2410.960 0.000 2414.500 1.120 ;
  LAYER metal1 ;
  RECT 2410.960 0.000 2414.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2402.280 0.000 2405.820 1.120 ;
  LAYER metal4 ;
  RECT 2402.280 0.000 2405.820 1.120 ;
  LAYER metal3 ;
  RECT 2402.280 0.000 2405.820 1.120 ;
  LAYER metal2 ;
  RECT 2402.280 0.000 2405.820 1.120 ;
  LAYER metal1 ;
  RECT 2402.280 0.000 2405.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2393.600 0.000 2397.140 1.120 ;
  LAYER metal4 ;
  RECT 2393.600 0.000 2397.140 1.120 ;
  LAYER metal3 ;
  RECT 2393.600 0.000 2397.140 1.120 ;
  LAYER metal2 ;
  RECT 2393.600 0.000 2397.140 1.120 ;
  LAYER metal1 ;
  RECT 2393.600 0.000 2397.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2384.920 0.000 2388.460 1.120 ;
  LAYER metal4 ;
  RECT 2384.920 0.000 2388.460 1.120 ;
  LAYER metal3 ;
  RECT 2384.920 0.000 2388.460 1.120 ;
  LAYER metal2 ;
  RECT 2384.920 0.000 2388.460 1.120 ;
  LAYER metal1 ;
  RECT 2384.920 0.000 2388.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2376.240 0.000 2379.780 1.120 ;
  LAYER metal4 ;
  RECT 2376.240 0.000 2379.780 1.120 ;
  LAYER metal3 ;
  RECT 2376.240 0.000 2379.780 1.120 ;
  LAYER metal2 ;
  RECT 2376.240 0.000 2379.780 1.120 ;
  LAYER metal1 ;
  RECT 2376.240 0.000 2379.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2323.540 0.000 2327.080 1.120 ;
  LAYER metal4 ;
  RECT 2323.540 0.000 2327.080 1.120 ;
  LAYER metal3 ;
  RECT 2323.540 0.000 2327.080 1.120 ;
  LAYER metal2 ;
  RECT 2323.540 0.000 2327.080 1.120 ;
  LAYER metal1 ;
  RECT 2323.540 0.000 2327.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2309.900 0.000 2313.440 1.120 ;
  LAYER metal4 ;
  RECT 2309.900 0.000 2313.440 1.120 ;
  LAYER metal3 ;
  RECT 2309.900 0.000 2313.440 1.120 ;
  LAYER metal2 ;
  RECT 2309.900 0.000 2313.440 1.120 ;
  LAYER metal1 ;
  RECT 2309.900 0.000 2313.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2295.640 0.000 2299.180 1.120 ;
  LAYER metal4 ;
  RECT 2295.640 0.000 2299.180 1.120 ;
  LAYER metal3 ;
  RECT 2295.640 0.000 2299.180 1.120 ;
  LAYER metal2 ;
  RECT 2295.640 0.000 2299.180 1.120 ;
  LAYER metal1 ;
  RECT 2295.640 0.000 2299.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2286.960 0.000 2290.500 1.120 ;
  LAYER metal4 ;
  RECT 2286.960 0.000 2290.500 1.120 ;
  LAYER metal3 ;
  RECT 2286.960 0.000 2290.500 1.120 ;
  LAYER metal2 ;
  RECT 2286.960 0.000 2290.500 1.120 ;
  LAYER metal1 ;
  RECT 2286.960 0.000 2290.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2278.280 0.000 2281.820 1.120 ;
  LAYER metal4 ;
  RECT 2278.280 0.000 2281.820 1.120 ;
  LAYER metal3 ;
  RECT 2278.280 0.000 2281.820 1.120 ;
  LAYER metal2 ;
  RECT 2278.280 0.000 2281.820 1.120 ;
  LAYER metal1 ;
  RECT 2278.280 0.000 2281.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2269.600 0.000 2273.140 1.120 ;
  LAYER metal4 ;
  RECT 2269.600 0.000 2273.140 1.120 ;
  LAYER metal3 ;
  RECT 2269.600 0.000 2273.140 1.120 ;
  LAYER metal2 ;
  RECT 2269.600 0.000 2273.140 1.120 ;
  LAYER metal1 ;
  RECT 2269.600 0.000 2273.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2226.200 0.000 2229.740 1.120 ;
  LAYER metal4 ;
  RECT 2226.200 0.000 2229.740 1.120 ;
  LAYER metal3 ;
  RECT 2226.200 0.000 2229.740 1.120 ;
  LAYER metal2 ;
  RECT 2226.200 0.000 2229.740 1.120 ;
  LAYER metal1 ;
  RECT 2226.200 0.000 2229.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2217.520 0.000 2221.060 1.120 ;
  LAYER metal4 ;
  RECT 2217.520 0.000 2221.060 1.120 ;
  LAYER metal3 ;
  RECT 2217.520 0.000 2221.060 1.120 ;
  LAYER metal2 ;
  RECT 2217.520 0.000 2221.060 1.120 ;
  LAYER metal1 ;
  RECT 2217.520 0.000 2221.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2208.840 0.000 2212.380 1.120 ;
  LAYER metal4 ;
  RECT 2208.840 0.000 2212.380 1.120 ;
  LAYER metal3 ;
  RECT 2208.840 0.000 2212.380 1.120 ;
  LAYER metal2 ;
  RECT 2208.840 0.000 2212.380 1.120 ;
  LAYER metal1 ;
  RECT 2208.840 0.000 2212.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2200.160 0.000 2203.700 1.120 ;
  LAYER metal4 ;
  RECT 2200.160 0.000 2203.700 1.120 ;
  LAYER metal3 ;
  RECT 2200.160 0.000 2203.700 1.120 ;
  LAYER metal2 ;
  RECT 2200.160 0.000 2203.700 1.120 ;
  LAYER metal1 ;
  RECT 2200.160 0.000 2203.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2191.480 0.000 2195.020 1.120 ;
  LAYER metal4 ;
  RECT 2191.480 0.000 2195.020 1.120 ;
  LAYER metal3 ;
  RECT 2191.480 0.000 2195.020 1.120 ;
  LAYER metal2 ;
  RECT 2191.480 0.000 2195.020 1.120 ;
  LAYER metal1 ;
  RECT 2191.480 0.000 2195.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2182.800 0.000 2186.340 1.120 ;
  LAYER metal4 ;
  RECT 2182.800 0.000 2186.340 1.120 ;
  LAYER metal3 ;
  RECT 2182.800 0.000 2186.340 1.120 ;
  LAYER metal2 ;
  RECT 2182.800 0.000 2186.340 1.120 ;
  LAYER metal1 ;
  RECT 2182.800 0.000 2186.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2139.400 0.000 2142.940 1.120 ;
  LAYER metal4 ;
  RECT 2139.400 0.000 2142.940 1.120 ;
  LAYER metal3 ;
  RECT 2139.400 0.000 2142.940 1.120 ;
  LAYER metal2 ;
  RECT 2139.400 0.000 2142.940 1.120 ;
  LAYER metal1 ;
  RECT 2139.400 0.000 2142.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2130.720 0.000 2134.260 1.120 ;
  LAYER metal4 ;
  RECT 2130.720 0.000 2134.260 1.120 ;
  LAYER metal3 ;
  RECT 2130.720 0.000 2134.260 1.120 ;
  LAYER metal2 ;
  RECT 2130.720 0.000 2134.260 1.120 ;
  LAYER metal1 ;
  RECT 2130.720 0.000 2134.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2122.040 0.000 2125.580 1.120 ;
  LAYER metal4 ;
  RECT 2122.040 0.000 2125.580 1.120 ;
  LAYER metal3 ;
  RECT 2122.040 0.000 2125.580 1.120 ;
  LAYER metal2 ;
  RECT 2122.040 0.000 2125.580 1.120 ;
  LAYER metal1 ;
  RECT 2122.040 0.000 2125.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2113.360 0.000 2116.900 1.120 ;
  LAYER metal4 ;
  RECT 2113.360 0.000 2116.900 1.120 ;
  LAYER metal3 ;
  RECT 2113.360 0.000 2116.900 1.120 ;
  LAYER metal2 ;
  RECT 2113.360 0.000 2116.900 1.120 ;
  LAYER metal1 ;
  RECT 2113.360 0.000 2116.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2104.680 0.000 2108.220 1.120 ;
  LAYER metal4 ;
  RECT 2104.680 0.000 2108.220 1.120 ;
  LAYER metal3 ;
  RECT 2104.680 0.000 2108.220 1.120 ;
  LAYER metal2 ;
  RECT 2104.680 0.000 2108.220 1.120 ;
  LAYER metal1 ;
  RECT 2104.680 0.000 2108.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2096.000 0.000 2099.540 1.120 ;
  LAYER metal4 ;
  RECT 2096.000 0.000 2099.540 1.120 ;
  LAYER metal3 ;
  RECT 2096.000 0.000 2099.540 1.120 ;
  LAYER metal2 ;
  RECT 2096.000 0.000 2099.540 1.120 ;
  LAYER metal1 ;
  RECT 2096.000 0.000 2099.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2052.600 0.000 2056.140 1.120 ;
  LAYER metal4 ;
  RECT 2052.600 0.000 2056.140 1.120 ;
  LAYER metal3 ;
  RECT 2052.600 0.000 2056.140 1.120 ;
  LAYER metal2 ;
  RECT 2052.600 0.000 2056.140 1.120 ;
  LAYER metal1 ;
  RECT 2052.600 0.000 2056.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2043.920 0.000 2047.460 1.120 ;
  LAYER metal4 ;
  RECT 2043.920 0.000 2047.460 1.120 ;
  LAYER metal3 ;
  RECT 2043.920 0.000 2047.460 1.120 ;
  LAYER metal2 ;
  RECT 2043.920 0.000 2047.460 1.120 ;
  LAYER metal1 ;
  RECT 2043.920 0.000 2047.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2035.240 0.000 2038.780 1.120 ;
  LAYER metal4 ;
  RECT 2035.240 0.000 2038.780 1.120 ;
  LAYER metal3 ;
  RECT 2035.240 0.000 2038.780 1.120 ;
  LAYER metal2 ;
  RECT 2035.240 0.000 2038.780 1.120 ;
  LAYER metal1 ;
  RECT 2035.240 0.000 2038.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2026.560 0.000 2030.100 1.120 ;
  LAYER metal4 ;
  RECT 2026.560 0.000 2030.100 1.120 ;
  LAYER metal3 ;
  RECT 2026.560 0.000 2030.100 1.120 ;
  LAYER metal2 ;
  RECT 2026.560 0.000 2030.100 1.120 ;
  LAYER metal1 ;
  RECT 2026.560 0.000 2030.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2017.880 0.000 2021.420 1.120 ;
  LAYER metal4 ;
  RECT 2017.880 0.000 2021.420 1.120 ;
  LAYER metal3 ;
  RECT 2017.880 0.000 2021.420 1.120 ;
  LAYER metal2 ;
  RECT 2017.880 0.000 2021.420 1.120 ;
  LAYER metal1 ;
  RECT 2017.880 0.000 2021.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2009.200 0.000 2012.740 1.120 ;
  LAYER metal4 ;
  RECT 2009.200 0.000 2012.740 1.120 ;
  LAYER metal3 ;
  RECT 2009.200 0.000 2012.740 1.120 ;
  LAYER metal2 ;
  RECT 2009.200 0.000 2012.740 1.120 ;
  LAYER metal1 ;
  RECT 2009.200 0.000 2012.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1965.800 0.000 1969.340 1.120 ;
  LAYER metal4 ;
  RECT 1965.800 0.000 1969.340 1.120 ;
  LAYER metal3 ;
  RECT 1965.800 0.000 1969.340 1.120 ;
  LAYER metal2 ;
  RECT 1965.800 0.000 1969.340 1.120 ;
  LAYER metal1 ;
  RECT 1965.800 0.000 1969.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1957.120 0.000 1960.660 1.120 ;
  LAYER metal4 ;
  RECT 1957.120 0.000 1960.660 1.120 ;
  LAYER metal3 ;
  RECT 1957.120 0.000 1960.660 1.120 ;
  LAYER metal2 ;
  RECT 1957.120 0.000 1960.660 1.120 ;
  LAYER metal1 ;
  RECT 1957.120 0.000 1960.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1948.440 0.000 1951.980 1.120 ;
  LAYER metal4 ;
  RECT 1948.440 0.000 1951.980 1.120 ;
  LAYER metal3 ;
  RECT 1948.440 0.000 1951.980 1.120 ;
  LAYER metal2 ;
  RECT 1948.440 0.000 1951.980 1.120 ;
  LAYER metal1 ;
  RECT 1948.440 0.000 1951.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1939.760 0.000 1943.300 1.120 ;
  LAYER metal4 ;
  RECT 1939.760 0.000 1943.300 1.120 ;
  LAYER metal3 ;
  RECT 1939.760 0.000 1943.300 1.120 ;
  LAYER metal2 ;
  RECT 1939.760 0.000 1943.300 1.120 ;
  LAYER metal1 ;
  RECT 1939.760 0.000 1943.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1931.080 0.000 1934.620 1.120 ;
  LAYER metal4 ;
  RECT 1931.080 0.000 1934.620 1.120 ;
  LAYER metal3 ;
  RECT 1931.080 0.000 1934.620 1.120 ;
  LAYER metal2 ;
  RECT 1931.080 0.000 1934.620 1.120 ;
  LAYER metal1 ;
  RECT 1931.080 0.000 1934.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1922.400 0.000 1925.940 1.120 ;
  LAYER metal4 ;
  RECT 1922.400 0.000 1925.940 1.120 ;
  LAYER metal3 ;
  RECT 1922.400 0.000 1925.940 1.120 ;
  LAYER metal2 ;
  RECT 1922.400 0.000 1925.940 1.120 ;
  LAYER metal1 ;
  RECT 1922.400 0.000 1925.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1859.160 0.000 1862.700 1.120 ;
  LAYER metal4 ;
  RECT 1859.160 0.000 1862.700 1.120 ;
  LAYER metal3 ;
  RECT 1859.160 0.000 1862.700 1.120 ;
  LAYER metal2 ;
  RECT 1859.160 0.000 1862.700 1.120 ;
  LAYER metal1 ;
  RECT 1859.160 0.000 1862.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1850.480 0.000 1854.020 1.120 ;
  LAYER metal4 ;
  RECT 1850.480 0.000 1854.020 1.120 ;
  LAYER metal3 ;
  RECT 1850.480 0.000 1854.020 1.120 ;
  LAYER metal2 ;
  RECT 1850.480 0.000 1854.020 1.120 ;
  LAYER metal1 ;
  RECT 1850.480 0.000 1854.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1793.440 0.000 1796.980 1.120 ;
  LAYER metal4 ;
  RECT 1793.440 0.000 1796.980 1.120 ;
  LAYER metal3 ;
  RECT 1793.440 0.000 1796.980 1.120 ;
  LAYER metal2 ;
  RECT 1793.440 0.000 1796.980 1.120 ;
  LAYER metal1 ;
  RECT 1793.440 0.000 1796.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1768.640 0.000 1772.180 1.120 ;
  LAYER metal4 ;
  RECT 1768.640 0.000 1772.180 1.120 ;
  LAYER metal3 ;
  RECT 1768.640 0.000 1772.180 1.120 ;
  LAYER metal2 ;
  RECT 1768.640 0.000 1772.180 1.120 ;
  LAYER metal1 ;
  RECT 1768.640 0.000 1772.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1742.600 0.000 1746.140 1.120 ;
  LAYER metal4 ;
  RECT 1742.600 0.000 1746.140 1.120 ;
  LAYER metal3 ;
  RECT 1742.600 0.000 1746.140 1.120 ;
  LAYER metal2 ;
  RECT 1742.600 0.000 1746.140 1.120 ;
  LAYER metal1 ;
  RECT 1742.600 0.000 1746.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1733.920 0.000 1737.460 1.120 ;
  LAYER metal4 ;
  RECT 1733.920 0.000 1737.460 1.120 ;
  LAYER metal3 ;
  RECT 1733.920 0.000 1737.460 1.120 ;
  LAYER metal2 ;
  RECT 1733.920 0.000 1737.460 1.120 ;
  LAYER metal1 ;
  RECT 1733.920 0.000 1737.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1690.520 0.000 1694.060 1.120 ;
  LAYER metal4 ;
  RECT 1690.520 0.000 1694.060 1.120 ;
  LAYER metal3 ;
  RECT 1690.520 0.000 1694.060 1.120 ;
  LAYER metal2 ;
  RECT 1690.520 0.000 1694.060 1.120 ;
  LAYER metal1 ;
  RECT 1690.520 0.000 1694.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1681.840 0.000 1685.380 1.120 ;
  LAYER metal4 ;
  RECT 1681.840 0.000 1685.380 1.120 ;
  LAYER metal3 ;
  RECT 1681.840 0.000 1685.380 1.120 ;
  LAYER metal2 ;
  RECT 1681.840 0.000 1685.380 1.120 ;
  LAYER metal1 ;
  RECT 1681.840 0.000 1685.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1673.160 0.000 1676.700 1.120 ;
  LAYER metal4 ;
  RECT 1673.160 0.000 1676.700 1.120 ;
  LAYER metal3 ;
  RECT 1673.160 0.000 1676.700 1.120 ;
  LAYER metal2 ;
  RECT 1673.160 0.000 1676.700 1.120 ;
  LAYER metal1 ;
  RECT 1673.160 0.000 1676.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1664.480 0.000 1668.020 1.120 ;
  LAYER metal4 ;
  RECT 1664.480 0.000 1668.020 1.120 ;
  LAYER metal3 ;
  RECT 1664.480 0.000 1668.020 1.120 ;
  LAYER metal2 ;
  RECT 1664.480 0.000 1668.020 1.120 ;
  LAYER metal1 ;
  RECT 1664.480 0.000 1668.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1655.800 0.000 1659.340 1.120 ;
  LAYER metal4 ;
  RECT 1655.800 0.000 1659.340 1.120 ;
  LAYER metal3 ;
  RECT 1655.800 0.000 1659.340 1.120 ;
  LAYER metal2 ;
  RECT 1655.800 0.000 1659.340 1.120 ;
  LAYER metal1 ;
  RECT 1655.800 0.000 1659.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1647.120 0.000 1650.660 1.120 ;
  LAYER metal4 ;
  RECT 1647.120 0.000 1650.660 1.120 ;
  LAYER metal3 ;
  RECT 1647.120 0.000 1650.660 1.120 ;
  LAYER metal2 ;
  RECT 1647.120 0.000 1650.660 1.120 ;
  LAYER metal1 ;
  RECT 1647.120 0.000 1650.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1603.720 0.000 1607.260 1.120 ;
  LAYER metal4 ;
  RECT 1603.720 0.000 1607.260 1.120 ;
  LAYER metal3 ;
  RECT 1603.720 0.000 1607.260 1.120 ;
  LAYER metal2 ;
  RECT 1603.720 0.000 1607.260 1.120 ;
  LAYER metal1 ;
  RECT 1603.720 0.000 1607.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1595.040 0.000 1598.580 1.120 ;
  LAYER metal4 ;
  RECT 1595.040 0.000 1598.580 1.120 ;
  LAYER metal3 ;
  RECT 1595.040 0.000 1598.580 1.120 ;
  LAYER metal2 ;
  RECT 1595.040 0.000 1598.580 1.120 ;
  LAYER metal1 ;
  RECT 1595.040 0.000 1598.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1586.360 0.000 1589.900 1.120 ;
  LAYER metal4 ;
  RECT 1586.360 0.000 1589.900 1.120 ;
  LAYER metal3 ;
  RECT 1586.360 0.000 1589.900 1.120 ;
  LAYER metal2 ;
  RECT 1586.360 0.000 1589.900 1.120 ;
  LAYER metal1 ;
  RECT 1586.360 0.000 1589.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1577.680 0.000 1581.220 1.120 ;
  LAYER metal4 ;
  RECT 1577.680 0.000 1581.220 1.120 ;
  LAYER metal3 ;
  RECT 1577.680 0.000 1581.220 1.120 ;
  LAYER metal2 ;
  RECT 1577.680 0.000 1581.220 1.120 ;
  LAYER metal1 ;
  RECT 1577.680 0.000 1581.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1569.000 0.000 1572.540 1.120 ;
  LAYER metal4 ;
  RECT 1569.000 0.000 1572.540 1.120 ;
  LAYER metal3 ;
  RECT 1569.000 0.000 1572.540 1.120 ;
  LAYER metal2 ;
  RECT 1569.000 0.000 1572.540 1.120 ;
  LAYER metal1 ;
  RECT 1569.000 0.000 1572.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1560.320 0.000 1563.860 1.120 ;
  LAYER metal4 ;
  RECT 1560.320 0.000 1563.860 1.120 ;
  LAYER metal3 ;
  RECT 1560.320 0.000 1563.860 1.120 ;
  LAYER metal2 ;
  RECT 1560.320 0.000 1563.860 1.120 ;
  LAYER metal1 ;
  RECT 1560.320 0.000 1563.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1516.920 0.000 1520.460 1.120 ;
  LAYER metal4 ;
  RECT 1516.920 0.000 1520.460 1.120 ;
  LAYER metal3 ;
  RECT 1516.920 0.000 1520.460 1.120 ;
  LAYER metal2 ;
  RECT 1516.920 0.000 1520.460 1.120 ;
  LAYER metal1 ;
  RECT 1516.920 0.000 1520.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1508.240 0.000 1511.780 1.120 ;
  LAYER metal4 ;
  RECT 1508.240 0.000 1511.780 1.120 ;
  LAYER metal3 ;
  RECT 1508.240 0.000 1511.780 1.120 ;
  LAYER metal2 ;
  RECT 1508.240 0.000 1511.780 1.120 ;
  LAYER metal1 ;
  RECT 1508.240 0.000 1511.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1499.560 0.000 1503.100 1.120 ;
  LAYER metal4 ;
  RECT 1499.560 0.000 1503.100 1.120 ;
  LAYER metal3 ;
  RECT 1499.560 0.000 1503.100 1.120 ;
  LAYER metal2 ;
  RECT 1499.560 0.000 1503.100 1.120 ;
  LAYER metal1 ;
  RECT 1499.560 0.000 1503.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1490.880 0.000 1494.420 1.120 ;
  LAYER metal4 ;
  RECT 1490.880 0.000 1494.420 1.120 ;
  LAYER metal3 ;
  RECT 1490.880 0.000 1494.420 1.120 ;
  LAYER metal2 ;
  RECT 1490.880 0.000 1494.420 1.120 ;
  LAYER metal1 ;
  RECT 1490.880 0.000 1494.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1482.200 0.000 1485.740 1.120 ;
  LAYER metal4 ;
  RECT 1482.200 0.000 1485.740 1.120 ;
  LAYER metal3 ;
  RECT 1482.200 0.000 1485.740 1.120 ;
  LAYER metal2 ;
  RECT 1482.200 0.000 1485.740 1.120 ;
  LAYER metal1 ;
  RECT 1482.200 0.000 1485.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1473.520 0.000 1477.060 1.120 ;
  LAYER metal4 ;
  RECT 1473.520 0.000 1477.060 1.120 ;
  LAYER metal3 ;
  RECT 1473.520 0.000 1477.060 1.120 ;
  LAYER metal2 ;
  RECT 1473.520 0.000 1477.060 1.120 ;
  LAYER metal1 ;
  RECT 1473.520 0.000 1477.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1430.120 0.000 1433.660 1.120 ;
  LAYER metal4 ;
  RECT 1430.120 0.000 1433.660 1.120 ;
  LAYER metal3 ;
  RECT 1430.120 0.000 1433.660 1.120 ;
  LAYER metal2 ;
  RECT 1430.120 0.000 1433.660 1.120 ;
  LAYER metal1 ;
  RECT 1430.120 0.000 1433.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1421.440 0.000 1424.980 1.120 ;
  LAYER metal4 ;
  RECT 1421.440 0.000 1424.980 1.120 ;
  LAYER metal3 ;
  RECT 1421.440 0.000 1424.980 1.120 ;
  LAYER metal2 ;
  RECT 1421.440 0.000 1424.980 1.120 ;
  LAYER metal1 ;
  RECT 1421.440 0.000 1424.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1412.760 0.000 1416.300 1.120 ;
  LAYER metal4 ;
  RECT 1412.760 0.000 1416.300 1.120 ;
  LAYER metal3 ;
  RECT 1412.760 0.000 1416.300 1.120 ;
  LAYER metal2 ;
  RECT 1412.760 0.000 1416.300 1.120 ;
  LAYER metal1 ;
  RECT 1412.760 0.000 1416.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1404.080 0.000 1407.620 1.120 ;
  LAYER metal4 ;
  RECT 1404.080 0.000 1407.620 1.120 ;
  LAYER metal3 ;
  RECT 1404.080 0.000 1407.620 1.120 ;
  LAYER metal2 ;
  RECT 1404.080 0.000 1407.620 1.120 ;
  LAYER metal1 ;
  RECT 1404.080 0.000 1407.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1395.400 0.000 1398.940 1.120 ;
  LAYER metal4 ;
  RECT 1395.400 0.000 1398.940 1.120 ;
  LAYER metal3 ;
  RECT 1395.400 0.000 1398.940 1.120 ;
  LAYER metal2 ;
  RECT 1395.400 0.000 1398.940 1.120 ;
  LAYER metal1 ;
  RECT 1395.400 0.000 1398.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1386.720 0.000 1390.260 1.120 ;
  LAYER metal4 ;
  RECT 1386.720 0.000 1390.260 1.120 ;
  LAYER metal3 ;
  RECT 1386.720 0.000 1390.260 1.120 ;
  LAYER metal2 ;
  RECT 1386.720 0.000 1390.260 1.120 ;
  LAYER metal1 ;
  RECT 1386.720 0.000 1390.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1338.980 0.000 1342.520 1.120 ;
  LAYER metal4 ;
  RECT 1338.980 0.000 1342.520 1.120 ;
  LAYER metal3 ;
  RECT 1338.980 0.000 1342.520 1.120 ;
  LAYER metal2 ;
  RECT 1338.980 0.000 1342.520 1.120 ;
  LAYER metal1 ;
  RECT 1338.980 0.000 1342.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1325.340 0.000 1328.880 1.120 ;
  LAYER metal4 ;
  RECT 1325.340 0.000 1328.880 1.120 ;
  LAYER metal3 ;
  RECT 1325.340 0.000 1328.880 1.120 ;
  LAYER metal2 ;
  RECT 1325.340 0.000 1328.880 1.120 ;
  LAYER metal1 ;
  RECT 1325.340 0.000 1328.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1311.700 0.000 1315.240 1.120 ;
  LAYER metal4 ;
  RECT 1311.700 0.000 1315.240 1.120 ;
  LAYER metal3 ;
  RECT 1311.700 0.000 1315.240 1.120 ;
  LAYER metal2 ;
  RECT 1311.700 0.000 1315.240 1.120 ;
  LAYER metal1 ;
  RECT 1311.700 0.000 1315.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1297.440 0.000 1300.980 1.120 ;
  LAYER metal4 ;
  RECT 1297.440 0.000 1300.980 1.120 ;
  LAYER metal3 ;
  RECT 1297.440 0.000 1300.980 1.120 ;
  LAYER metal2 ;
  RECT 1297.440 0.000 1300.980 1.120 ;
  LAYER metal1 ;
  RECT 1297.440 0.000 1300.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1288.760 0.000 1292.300 1.120 ;
  LAYER metal4 ;
  RECT 1288.760 0.000 1292.300 1.120 ;
  LAYER metal3 ;
  RECT 1288.760 0.000 1292.300 1.120 ;
  LAYER metal2 ;
  RECT 1288.760 0.000 1292.300 1.120 ;
  LAYER metal1 ;
  RECT 1288.760 0.000 1292.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1280.080 0.000 1283.620 1.120 ;
  LAYER metal4 ;
  RECT 1280.080 0.000 1283.620 1.120 ;
  LAYER metal3 ;
  RECT 1280.080 0.000 1283.620 1.120 ;
  LAYER metal2 ;
  RECT 1280.080 0.000 1283.620 1.120 ;
  LAYER metal1 ;
  RECT 1280.080 0.000 1283.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1236.680 0.000 1240.220 1.120 ;
  LAYER metal4 ;
  RECT 1236.680 0.000 1240.220 1.120 ;
  LAYER metal3 ;
  RECT 1236.680 0.000 1240.220 1.120 ;
  LAYER metal2 ;
  RECT 1236.680 0.000 1240.220 1.120 ;
  LAYER metal1 ;
  RECT 1236.680 0.000 1240.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1228.000 0.000 1231.540 1.120 ;
  LAYER metal4 ;
  RECT 1228.000 0.000 1231.540 1.120 ;
  LAYER metal3 ;
  RECT 1228.000 0.000 1231.540 1.120 ;
  LAYER metal2 ;
  RECT 1228.000 0.000 1231.540 1.120 ;
  LAYER metal1 ;
  RECT 1228.000 0.000 1231.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1219.320 0.000 1222.860 1.120 ;
  LAYER metal4 ;
  RECT 1219.320 0.000 1222.860 1.120 ;
  LAYER metal3 ;
  RECT 1219.320 0.000 1222.860 1.120 ;
  LAYER metal2 ;
  RECT 1219.320 0.000 1222.860 1.120 ;
  LAYER metal1 ;
  RECT 1219.320 0.000 1222.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1210.640 0.000 1214.180 1.120 ;
  LAYER metal4 ;
  RECT 1210.640 0.000 1214.180 1.120 ;
  LAYER metal3 ;
  RECT 1210.640 0.000 1214.180 1.120 ;
  LAYER metal2 ;
  RECT 1210.640 0.000 1214.180 1.120 ;
  LAYER metal1 ;
  RECT 1210.640 0.000 1214.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1201.960 0.000 1205.500 1.120 ;
  LAYER metal4 ;
  RECT 1201.960 0.000 1205.500 1.120 ;
  LAYER metal3 ;
  RECT 1201.960 0.000 1205.500 1.120 ;
  LAYER metal2 ;
  RECT 1201.960 0.000 1205.500 1.120 ;
  LAYER metal1 ;
  RECT 1201.960 0.000 1205.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1193.280 0.000 1196.820 1.120 ;
  LAYER metal4 ;
  RECT 1193.280 0.000 1196.820 1.120 ;
  LAYER metal3 ;
  RECT 1193.280 0.000 1196.820 1.120 ;
  LAYER metal2 ;
  RECT 1193.280 0.000 1196.820 1.120 ;
  LAYER metal1 ;
  RECT 1193.280 0.000 1196.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1149.880 0.000 1153.420 1.120 ;
  LAYER metal4 ;
  RECT 1149.880 0.000 1153.420 1.120 ;
  LAYER metal3 ;
  RECT 1149.880 0.000 1153.420 1.120 ;
  LAYER metal2 ;
  RECT 1149.880 0.000 1153.420 1.120 ;
  LAYER metal1 ;
  RECT 1149.880 0.000 1153.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1141.200 0.000 1144.740 1.120 ;
  LAYER metal4 ;
  RECT 1141.200 0.000 1144.740 1.120 ;
  LAYER metal3 ;
  RECT 1141.200 0.000 1144.740 1.120 ;
  LAYER metal2 ;
  RECT 1141.200 0.000 1144.740 1.120 ;
  LAYER metal1 ;
  RECT 1141.200 0.000 1144.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1132.520 0.000 1136.060 1.120 ;
  LAYER metal4 ;
  RECT 1132.520 0.000 1136.060 1.120 ;
  LAYER metal3 ;
  RECT 1132.520 0.000 1136.060 1.120 ;
  LAYER metal2 ;
  RECT 1132.520 0.000 1136.060 1.120 ;
  LAYER metal1 ;
  RECT 1132.520 0.000 1136.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1123.840 0.000 1127.380 1.120 ;
  LAYER metal4 ;
  RECT 1123.840 0.000 1127.380 1.120 ;
  LAYER metal3 ;
  RECT 1123.840 0.000 1127.380 1.120 ;
  LAYER metal2 ;
  RECT 1123.840 0.000 1127.380 1.120 ;
  LAYER metal1 ;
  RECT 1123.840 0.000 1127.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1115.160 0.000 1118.700 1.120 ;
  LAYER metal4 ;
  RECT 1115.160 0.000 1118.700 1.120 ;
  LAYER metal3 ;
  RECT 1115.160 0.000 1118.700 1.120 ;
  LAYER metal2 ;
  RECT 1115.160 0.000 1118.700 1.120 ;
  LAYER metal1 ;
  RECT 1115.160 0.000 1118.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1106.480 0.000 1110.020 1.120 ;
  LAYER metal4 ;
  RECT 1106.480 0.000 1110.020 1.120 ;
  LAYER metal3 ;
  RECT 1106.480 0.000 1110.020 1.120 ;
  LAYER metal2 ;
  RECT 1106.480 0.000 1110.020 1.120 ;
  LAYER metal1 ;
  RECT 1106.480 0.000 1110.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1063.080 0.000 1066.620 1.120 ;
  LAYER metal4 ;
  RECT 1063.080 0.000 1066.620 1.120 ;
  LAYER metal3 ;
  RECT 1063.080 0.000 1066.620 1.120 ;
  LAYER metal2 ;
  RECT 1063.080 0.000 1066.620 1.120 ;
  LAYER metal1 ;
  RECT 1063.080 0.000 1066.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1054.400 0.000 1057.940 1.120 ;
  LAYER metal4 ;
  RECT 1054.400 0.000 1057.940 1.120 ;
  LAYER metal3 ;
  RECT 1054.400 0.000 1057.940 1.120 ;
  LAYER metal2 ;
  RECT 1054.400 0.000 1057.940 1.120 ;
  LAYER metal1 ;
  RECT 1054.400 0.000 1057.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1045.720 0.000 1049.260 1.120 ;
  LAYER metal4 ;
  RECT 1045.720 0.000 1049.260 1.120 ;
  LAYER metal3 ;
  RECT 1045.720 0.000 1049.260 1.120 ;
  LAYER metal2 ;
  RECT 1045.720 0.000 1049.260 1.120 ;
  LAYER metal1 ;
  RECT 1045.720 0.000 1049.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1037.040 0.000 1040.580 1.120 ;
  LAYER metal4 ;
  RECT 1037.040 0.000 1040.580 1.120 ;
  LAYER metal3 ;
  RECT 1037.040 0.000 1040.580 1.120 ;
  LAYER metal2 ;
  RECT 1037.040 0.000 1040.580 1.120 ;
  LAYER metal1 ;
  RECT 1037.040 0.000 1040.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1028.360 0.000 1031.900 1.120 ;
  LAYER metal4 ;
  RECT 1028.360 0.000 1031.900 1.120 ;
  LAYER metal3 ;
  RECT 1028.360 0.000 1031.900 1.120 ;
  LAYER metal2 ;
  RECT 1028.360 0.000 1031.900 1.120 ;
  LAYER metal1 ;
  RECT 1028.360 0.000 1031.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1019.680 0.000 1023.220 1.120 ;
  LAYER metal4 ;
  RECT 1019.680 0.000 1023.220 1.120 ;
  LAYER metal3 ;
  RECT 1019.680 0.000 1023.220 1.120 ;
  LAYER metal2 ;
  RECT 1019.680 0.000 1023.220 1.120 ;
  LAYER metal1 ;
  RECT 1019.680 0.000 1023.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 976.280 0.000 979.820 1.120 ;
  LAYER metal4 ;
  RECT 976.280 0.000 979.820 1.120 ;
  LAYER metal3 ;
  RECT 976.280 0.000 979.820 1.120 ;
  LAYER metal2 ;
  RECT 976.280 0.000 979.820 1.120 ;
  LAYER metal1 ;
  RECT 976.280 0.000 979.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 967.600 0.000 971.140 1.120 ;
  LAYER metal4 ;
  RECT 967.600 0.000 971.140 1.120 ;
  LAYER metal3 ;
  RECT 967.600 0.000 971.140 1.120 ;
  LAYER metal2 ;
  RECT 967.600 0.000 971.140 1.120 ;
  LAYER metal1 ;
  RECT 967.600 0.000 971.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 958.920 0.000 962.460 1.120 ;
  LAYER metal4 ;
  RECT 958.920 0.000 962.460 1.120 ;
  LAYER metal3 ;
  RECT 958.920 0.000 962.460 1.120 ;
  LAYER metal2 ;
  RECT 958.920 0.000 962.460 1.120 ;
  LAYER metal1 ;
  RECT 958.920 0.000 962.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 950.240 0.000 953.780 1.120 ;
  LAYER metal4 ;
  RECT 950.240 0.000 953.780 1.120 ;
  LAYER metal3 ;
  RECT 950.240 0.000 953.780 1.120 ;
  LAYER metal2 ;
  RECT 950.240 0.000 953.780 1.120 ;
  LAYER metal1 ;
  RECT 950.240 0.000 953.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 941.560 0.000 945.100 1.120 ;
  LAYER metal4 ;
  RECT 941.560 0.000 945.100 1.120 ;
  LAYER metal3 ;
  RECT 941.560 0.000 945.100 1.120 ;
  LAYER metal2 ;
  RECT 941.560 0.000 945.100 1.120 ;
  LAYER metal1 ;
  RECT 941.560 0.000 945.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 932.880 0.000 936.420 1.120 ;
  LAYER metal4 ;
  RECT 932.880 0.000 936.420 1.120 ;
  LAYER metal3 ;
  RECT 932.880 0.000 936.420 1.120 ;
  LAYER metal2 ;
  RECT 932.880 0.000 936.420 1.120 ;
  LAYER metal1 ;
  RECT 932.880 0.000 936.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 869.640 0.000 873.180 1.120 ;
  LAYER metal4 ;
  RECT 869.640 0.000 873.180 1.120 ;
  LAYER metal3 ;
  RECT 869.640 0.000 873.180 1.120 ;
  LAYER metal2 ;
  RECT 869.640 0.000 873.180 1.120 ;
  LAYER metal1 ;
  RECT 869.640 0.000 873.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 860.960 0.000 864.500 1.120 ;
  LAYER metal4 ;
  RECT 860.960 0.000 864.500 1.120 ;
  LAYER metal3 ;
  RECT 860.960 0.000 864.500 1.120 ;
  LAYER metal2 ;
  RECT 860.960 0.000 864.500 1.120 ;
  LAYER metal1 ;
  RECT 860.960 0.000 864.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 852.280 0.000 855.820 1.120 ;
  LAYER metal4 ;
  RECT 852.280 0.000 855.820 1.120 ;
  LAYER metal3 ;
  RECT 852.280 0.000 855.820 1.120 ;
  LAYER metal2 ;
  RECT 852.280 0.000 855.820 1.120 ;
  LAYER metal1 ;
  RECT 852.280 0.000 855.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 843.600 0.000 847.140 1.120 ;
  LAYER metal4 ;
  RECT 843.600 0.000 847.140 1.120 ;
  LAYER metal3 ;
  RECT 843.600 0.000 847.140 1.120 ;
  LAYER metal2 ;
  RECT 843.600 0.000 847.140 1.120 ;
  LAYER metal1 ;
  RECT 843.600 0.000 847.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 834.920 0.000 838.460 1.120 ;
  LAYER metal4 ;
  RECT 834.920 0.000 838.460 1.120 ;
  LAYER metal3 ;
  RECT 834.920 0.000 838.460 1.120 ;
  LAYER metal2 ;
  RECT 834.920 0.000 838.460 1.120 ;
  LAYER metal1 ;
  RECT 834.920 0.000 838.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 826.240 0.000 829.780 1.120 ;
  LAYER metal4 ;
  RECT 826.240 0.000 829.780 1.120 ;
  LAYER metal3 ;
  RECT 826.240 0.000 829.780 1.120 ;
  LAYER metal2 ;
  RECT 826.240 0.000 829.780 1.120 ;
  LAYER metal1 ;
  RECT 826.240 0.000 829.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 782.840 0.000 786.380 1.120 ;
  LAYER metal4 ;
  RECT 782.840 0.000 786.380 1.120 ;
  LAYER metal3 ;
  RECT 782.840 0.000 786.380 1.120 ;
  LAYER metal2 ;
  RECT 782.840 0.000 786.380 1.120 ;
  LAYER metal1 ;
  RECT 782.840 0.000 786.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 774.160 0.000 777.700 1.120 ;
  LAYER metal4 ;
  RECT 774.160 0.000 777.700 1.120 ;
  LAYER metal3 ;
  RECT 774.160 0.000 777.700 1.120 ;
  LAYER metal2 ;
  RECT 774.160 0.000 777.700 1.120 ;
  LAYER metal1 ;
  RECT 774.160 0.000 777.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 765.480 0.000 769.020 1.120 ;
  LAYER metal4 ;
  RECT 765.480 0.000 769.020 1.120 ;
  LAYER metal3 ;
  RECT 765.480 0.000 769.020 1.120 ;
  LAYER metal2 ;
  RECT 765.480 0.000 769.020 1.120 ;
  LAYER metal1 ;
  RECT 765.480 0.000 769.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 756.800 0.000 760.340 1.120 ;
  LAYER metal4 ;
  RECT 756.800 0.000 760.340 1.120 ;
  LAYER metal3 ;
  RECT 756.800 0.000 760.340 1.120 ;
  LAYER metal2 ;
  RECT 756.800 0.000 760.340 1.120 ;
  LAYER metal1 ;
  RECT 756.800 0.000 760.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 748.120 0.000 751.660 1.120 ;
  LAYER metal4 ;
  RECT 748.120 0.000 751.660 1.120 ;
  LAYER metal3 ;
  RECT 748.120 0.000 751.660 1.120 ;
  LAYER metal2 ;
  RECT 748.120 0.000 751.660 1.120 ;
  LAYER metal1 ;
  RECT 748.120 0.000 751.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 739.440 0.000 742.980 1.120 ;
  LAYER metal4 ;
  RECT 739.440 0.000 742.980 1.120 ;
  LAYER metal3 ;
  RECT 739.440 0.000 742.980 1.120 ;
  LAYER metal2 ;
  RECT 739.440 0.000 742.980 1.120 ;
  LAYER metal1 ;
  RECT 739.440 0.000 742.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 696.040 0.000 699.580 1.120 ;
  LAYER metal4 ;
  RECT 696.040 0.000 699.580 1.120 ;
  LAYER metal3 ;
  RECT 696.040 0.000 699.580 1.120 ;
  LAYER metal2 ;
  RECT 696.040 0.000 699.580 1.120 ;
  LAYER metal1 ;
  RECT 696.040 0.000 699.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 687.360 0.000 690.900 1.120 ;
  LAYER metal4 ;
  RECT 687.360 0.000 690.900 1.120 ;
  LAYER metal3 ;
  RECT 687.360 0.000 690.900 1.120 ;
  LAYER metal2 ;
  RECT 687.360 0.000 690.900 1.120 ;
  LAYER metal1 ;
  RECT 687.360 0.000 690.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 678.680 0.000 682.220 1.120 ;
  LAYER metal4 ;
  RECT 678.680 0.000 682.220 1.120 ;
  LAYER metal3 ;
  RECT 678.680 0.000 682.220 1.120 ;
  LAYER metal2 ;
  RECT 678.680 0.000 682.220 1.120 ;
  LAYER metal1 ;
  RECT 678.680 0.000 682.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 670.000 0.000 673.540 1.120 ;
  LAYER metal4 ;
  RECT 670.000 0.000 673.540 1.120 ;
  LAYER metal3 ;
  RECT 670.000 0.000 673.540 1.120 ;
  LAYER metal2 ;
  RECT 670.000 0.000 673.540 1.120 ;
  LAYER metal1 ;
  RECT 670.000 0.000 673.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 661.320 0.000 664.860 1.120 ;
  LAYER metal4 ;
  RECT 661.320 0.000 664.860 1.120 ;
  LAYER metal3 ;
  RECT 661.320 0.000 664.860 1.120 ;
  LAYER metal2 ;
  RECT 661.320 0.000 664.860 1.120 ;
  LAYER metal1 ;
  RECT 661.320 0.000 664.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 652.640 0.000 656.180 1.120 ;
  LAYER metal4 ;
  RECT 652.640 0.000 656.180 1.120 ;
  LAYER metal3 ;
  RECT 652.640 0.000 656.180 1.120 ;
  LAYER metal2 ;
  RECT 652.640 0.000 656.180 1.120 ;
  LAYER metal1 ;
  RECT 652.640 0.000 656.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 609.240 0.000 612.780 1.120 ;
  LAYER metal4 ;
  RECT 609.240 0.000 612.780 1.120 ;
  LAYER metal3 ;
  RECT 609.240 0.000 612.780 1.120 ;
  LAYER metal2 ;
  RECT 609.240 0.000 612.780 1.120 ;
  LAYER metal1 ;
  RECT 609.240 0.000 612.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 600.560 0.000 604.100 1.120 ;
  LAYER metal4 ;
  RECT 600.560 0.000 604.100 1.120 ;
  LAYER metal3 ;
  RECT 600.560 0.000 604.100 1.120 ;
  LAYER metal2 ;
  RECT 600.560 0.000 604.100 1.120 ;
  LAYER metal1 ;
  RECT 600.560 0.000 604.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 591.880 0.000 595.420 1.120 ;
  LAYER metal4 ;
  RECT 591.880 0.000 595.420 1.120 ;
  LAYER metal3 ;
  RECT 591.880 0.000 595.420 1.120 ;
  LAYER metal2 ;
  RECT 591.880 0.000 595.420 1.120 ;
  LAYER metal1 ;
  RECT 591.880 0.000 595.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 583.200 0.000 586.740 1.120 ;
  LAYER metal4 ;
  RECT 583.200 0.000 586.740 1.120 ;
  LAYER metal3 ;
  RECT 583.200 0.000 586.740 1.120 ;
  LAYER metal2 ;
  RECT 583.200 0.000 586.740 1.120 ;
  LAYER metal1 ;
  RECT 583.200 0.000 586.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 574.520 0.000 578.060 1.120 ;
  LAYER metal4 ;
  RECT 574.520 0.000 578.060 1.120 ;
  LAYER metal3 ;
  RECT 574.520 0.000 578.060 1.120 ;
  LAYER metal2 ;
  RECT 574.520 0.000 578.060 1.120 ;
  LAYER metal1 ;
  RECT 574.520 0.000 578.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER metal4 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER metal3 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER metal2 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER metal1 ;
  RECT 565.840 0.000 569.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 522.440 0.000 525.980 1.120 ;
  LAYER metal4 ;
  RECT 522.440 0.000 525.980 1.120 ;
  LAYER metal3 ;
  RECT 522.440 0.000 525.980 1.120 ;
  LAYER metal2 ;
  RECT 522.440 0.000 525.980 1.120 ;
  LAYER metal1 ;
  RECT 522.440 0.000 525.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 513.760 0.000 517.300 1.120 ;
  LAYER metal4 ;
  RECT 513.760 0.000 517.300 1.120 ;
  LAYER metal3 ;
  RECT 513.760 0.000 517.300 1.120 ;
  LAYER metal2 ;
  RECT 513.760 0.000 517.300 1.120 ;
  LAYER metal1 ;
  RECT 513.760 0.000 517.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 505.080 0.000 508.620 1.120 ;
  LAYER metal4 ;
  RECT 505.080 0.000 508.620 1.120 ;
  LAYER metal3 ;
  RECT 505.080 0.000 508.620 1.120 ;
  LAYER metal2 ;
  RECT 505.080 0.000 508.620 1.120 ;
  LAYER metal1 ;
  RECT 505.080 0.000 508.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 496.400 0.000 499.940 1.120 ;
  LAYER metal4 ;
  RECT 496.400 0.000 499.940 1.120 ;
  LAYER metal3 ;
  RECT 496.400 0.000 499.940 1.120 ;
  LAYER metal2 ;
  RECT 496.400 0.000 499.940 1.120 ;
  LAYER metal1 ;
  RECT 496.400 0.000 499.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 487.720 0.000 491.260 1.120 ;
  LAYER metal4 ;
  RECT 487.720 0.000 491.260 1.120 ;
  LAYER metal3 ;
  RECT 487.720 0.000 491.260 1.120 ;
  LAYER metal2 ;
  RECT 487.720 0.000 491.260 1.120 ;
  LAYER metal1 ;
  RECT 487.720 0.000 491.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 474.080 0.000 477.620 1.120 ;
  LAYER metal4 ;
  RECT 474.080 0.000 477.620 1.120 ;
  LAYER metal3 ;
  RECT 474.080 0.000 477.620 1.120 ;
  LAYER metal2 ;
  RECT 474.080 0.000 477.620 1.120 ;
  LAYER metal1 ;
  RECT 474.080 0.000 477.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 415.180 0.000 418.720 1.120 ;
  LAYER metal4 ;
  RECT 415.180 0.000 418.720 1.120 ;
  LAYER metal3 ;
  RECT 415.180 0.000 418.720 1.120 ;
  LAYER metal2 ;
  RECT 415.180 0.000 418.720 1.120 ;
  LAYER metal1 ;
  RECT 415.180 0.000 418.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 406.500 0.000 410.040 1.120 ;
  LAYER metal4 ;
  RECT 406.500 0.000 410.040 1.120 ;
  LAYER metal3 ;
  RECT 406.500 0.000 410.040 1.120 ;
  LAYER metal2 ;
  RECT 406.500 0.000 410.040 1.120 ;
  LAYER metal1 ;
  RECT 406.500 0.000 410.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 397.820 0.000 401.360 1.120 ;
  LAYER metal4 ;
  RECT 397.820 0.000 401.360 1.120 ;
  LAYER metal3 ;
  RECT 397.820 0.000 401.360 1.120 ;
  LAYER metal2 ;
  RECT 397.820 0.000 401.360 1.120 ;
  LAYER metal1 ;
  RECT 397.820 0.000 401.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 389.140 0.000 392.680 1.120 ;
  LAYER metal4 ;
  RECT 389.140 0.000 392.680 1.120 ;
  LAYER metal3 ;
  RECT 389.140 0.000 392.680 1.120 ;
  LAYER metal2 ;
  RECT 389.140 0.000 392.680 1.120 ;
  LAYER metal1 ;
  RECT 389.140 0.000 392.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 380.460 0.000 384.000 1.120 ;
  LAYER metal4 ;
  RECT 380.460 0.000 384.000 1.120 ;
  LAYER metal3 ;
  RECT 380.460 0.000 384.000 1.120 ;
  LAYER metal2 ;
  RECT 380.460 0.000 384.000 1.120 ;
  LAYER metal1 ;
  RECT 380.460 0.000 384.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 371.780 0.000 375.320 1.120 ;
  LAYER metal4 ;
  RECT 371.780 0.000 375.320 1.120 ;
  LAYER metal3 ;
  RECT 371.780 0.000 375.320 1.120 ;
  LAYER metal2 ;
  RECT 371.780 0.000 375.320 1.120 ;
  LAYER metal1 ;
  RECT 371.780 0.000 375.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER metal4 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER metal3 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER metal2 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER metal1 ;
  RECT 328.380 0.000 331.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 319.700 0.000 323.240 1.120 ;
  LAYER metal4 ;
  RECT 319.700 0.000 323.240 1.120 ;
  LAYER metal3 ;
  RECT 319.700 0.000 323.240 1.120 ;
  LAYER metal2 ;
  RECT 319.700 0.000 323.240 1.120 ;
  LAYER metal1 ;
  RECT 319.700 0.000 323.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 311.020 0.000 314.560 1.120 ;
  LAYER metal4 ;
  RECT 311.020 0.000 314.560 1.120 ;
  LAYER metal3 ;
  RECT 311.020 0.000 314.560 1.120 ;
  LAYER metal2 ;
  RECT 311.020 0.000 314.560 1.120 ;
  LAYER metal1 ;
  RECT 311.020 0.000 314.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 302.340 0.000 305.880 1.120 ;
  LAYER metal4 ;
  RECT 302.340 0.000 305.880 1.120 ;
  LAYER metal3 ;
  RECT 302.340 0.000 305.880 1.120 ;
  LAYER metal2 ;
  RECT 302.340 0.000 305.880 1.120 ;
  LAYER metal1 ;
  RECT 302.340 0.000 305.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 293.660 0.000 297.200 1.120 ;
  LAYER metal4 ;
  RECT 293.660 0.000 297.200 1.120 ;
  LAYER metal3 ;
  RECT 293.660 0.000 297.200 1.120 ;
  LAYER metal2 ;
  RECT 293.660 0.000 297.200 1.120 ;
  LAYER metal1 ;
  RECT 293.660 0.000 297.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 284.980 0.000 288.520 1.120 ;
  LAYER metal4 ;
  RECT 284.980 0.000 288.520 1.120 ;
  LAYER metal3 ;
  RECT 284.980 0.000 288.520 1.120 ;
  LAYER metal2 ;
  RECT 284.980 0.000 288.520 1.120 ;
  LAYER metal1 ;
  RECT 284.980 0.000 288.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 241.580 0.000 245.120 1.120 ;
  LAYER metal4 ;
  RECT 241.580 0.000 245.120 1.120 ;
  LAYER metal3 ;
  RECT 241.580 0.000 245.120 1.120 ;
  LAYER metal2 ;
  RECT 241.580 0.000 245.120 1.120 ;
  LAYER metal1 ;
  RECT 241.580 0.000 245.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 232.900 0.000 236.440 1.120 ;
  LAYER metal4 ;
  RECT 232.900 0.000 236.440 1.120 ;
  LAYER metal3 ;
  RECT 232.900 0.000 236.440 1.120 ;
  LAYER metal2 ;
  RECT 232.900 0.000 236.440 1.120 ;
  LAYER metal1 ;
  RECT 232.900 0.000 236.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 224.220 0.000 227.760 1.120 ;
  LAYER metal4 ;
  RECT 224.220 0.000 227.760 1.120 ;
  LAYER metal3 ;
  RECT 224.220 0.000 227.760 1.120 ;
  LAYER metal2 ;
  RECT 224.220 0.000 227.760 1.120 ;
  LAYER metal1 ;
  RECT 224.220 0.000 227.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 215.540 0.000 219.080 1.120 ;
  LAYER metal4 ;
  RECT 215.540 0.000 219.080 1.120 ;
  LAYER metal3 ;
  RECT 215.540 0.000 219.080 1.120 ;
  LAYER metal2 ;
  RECT 215.540 0.000 219.080 1.120 ;
  LAYER metal1 ;
  RECT 215.540 0.000 219.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 206.860 0.000 210.400 1.120 ;
  LAYER metal4 ;
  RECT 206.860 0.000 210.400 1.120 ;
  LAYER metal3 ;
  RECT 206.860 0.000 210.400 1.120 ;
  LAYER metal2 ;
  RECT 206.860 0.000 210.400 1.120 ;
  LAYER metal1 ;
  RECT 206.860 0.000 210.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 198.180 0.000 201.720 1.120 ;
  LAYER metal4 ;
  RECT 198.180 0.000 201.720 1.120 ;
  LAYER metal3 ;
  RECT 198.180 0.000 201.720 1.120 ;
  LAYER metal2 ;
  RECT 198.180 0.000 201.720 1.120 ;
  LAYER metal1 ;
  RECT 198.180 0.000 201.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 154.780 0.000 158.320 1.120 ;
  LAYER metal4 ;
  RECT 154.780 0.000 158.320 1.120 ;
  LAYER metal3 ;
  RECT 154.780 0.000 158.320 1.120 ;
  LAYER metal2 ;
  RECT 154.780 0.000 158.320 1.120 ;
  LAYER metal1 ;
  RECT 154.780 0.000 158.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 146.100 0.000 149.640 1.120 ;
  LAYER metal4 ;
  RECT 146.100 0.000 149.640 1.120 ;
  LAYER metal3 ;
  RECT 146.100 0.000 149.640 1.120 ;
  LAYER metal2 ;
  RECT 146.100 0.000 149.640 1.120 ;
  LAYER metal1 ;
  RECT 146.100 0.000 149.640 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 137.420 0.000 140.960 1.120 ;
  LAYER metal4 ;
  RECT 137.420 0.000 140.960 1.120 ;
  LAYER metal3 ;
  RECT 137.420 0.000 140.960 1.120 ;
  LAYER metal2 ;
  RECT 137.420 0.000 140.960 1.120 ;
  LAYER metal1 ;
  RECT 137.420 0.000 140.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 128.740 0.000 132.280 1.120 ;
  LAYER metal4 ;
  RECT 128.740 0.000 132.280 1.120 ;
  LAYER metal3 ;
  RECT 128.740 0.000 132.280 1.120 ;
  LAYER metal2 ;
  RECT 128.740 0.000 132.280 1.120 ;
  LAYER metal1 ;
  RECT 128.740 0.000 132.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 120.060 0.000 123.600 1.120 ;
  LAYER metal4 ;
  RECT 120.060 0.000 123.600 1.120 ;
  LAYER metal3 ;
  RECT 120.060 0.000 123.600 1.120 ;
  LAYER metal2 ;
  RECT 120.060 0.000 123.600 1.120 ;
  LAYER metal1 ;
  RECT 120.060 0.000 123.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 111.380 0.000 114.920 1.120 ;
  LAYER metal4 ;
  RECT 111.380 0.000 114.920 1.120 ;
  LAYER metal3 ;
  RECT 111.380 0.000 114.920 1.120 ;
  LAYER metal2 ;
  RECT 111.380 0.000 114.920 1.120 ;
  LAYER metal1 ;
  RECT 111.380 0.000 114.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 67.980 0.000 71.520 1.120 ;
  LAYER metal4 ;
  RECT 67.980 0.000 71.520 1.120 ;
  LAYER metal3 ;
  RECT 67.980 0.000 71.520 1.120 ;
  LAYER metal2 ;
  RECT 67.980 0.000 71.520 1.120 ;
  LAYER metal1 ;
  RECT 67.980 0.000 71.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER metal4 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER metal3 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER metal2 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER metal1 ;
  RECT 59.300 0.000 62.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER metal4 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER metal3 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER metal2 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER metal1 ;
  RECT 46.280 0.000 49.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER metal4 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER metal3 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER metal2 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER metal1 ;
  RECT 32.640 0.000 36.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 19.000 0.000 22.540 1.120 ;
  LAYER metal4 ;
  RECT 19.000 0.000 22.540 1.120 ;
  LAYER metal3 ;
  RECT 19.000 0.000 22.540 1.120 ;
  LAYER metal2 ;
  RECT 19.000 0.000 22.540 1.120 ;
  LAYER metal1 ;
  RECT 19.000 0.000 22.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER metal4 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER metal3 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER metal2 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER metal1 ;
  RECT 7.220 0.000 10.760 1.120 ;
 END
END VCC
PIN DIB15
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3212.280 1710.800 3213.400 1711.920 ;
  LAYER metal4 ;
  RECT 3212.280 1710.800 3213.400 1711.920 ;
  LAYER metal3 ;
  RECT 3212.280 1710.800 3213.400 1711.920 ;
  LAYER metal2 ;
  RECT 3212.280 1710.800 3213.400 1711.920 ;
  LAYER metal1 ;
  RECT 3212.280 1710.800 3213.400 1711.920 ;
 END
END DIB15
PIN DOB15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3199.260 1710.800 3200.380 1711.920 ;
  LAYER metal4 ;
  RECT 3199.260 1710.800 3200.380 1711.920 ;
  LAYER metal3 ;
  RECT 3199.260 1710.800 3200.380 1711.920 ;
  LAYER metal2 ;
  RECT 3199.260 1710.800 3200.380 1711.920 ;
  LAYER metal1 ;
  RECT 3199.260 1710.800 3200.380 1711.920 ;
 END
END DOB15
PIN DIB14
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3185.620 1710.800 3186.740 1711.920 ;
  LAYER metal4 ;
  RECT 3185.620 1710.800 3186.740 1711.920 ;
  LAYER metal3 ;
  RECT 3185.620 1710.800 3186.740 1711.920 ;
  LAYER metal2 ;
  RECT 3185.620 1710.800 3186.740 1711.920 ;
  LAYER metal1 ;
  RECT 3185.620 1710.800 3186.740 1711.920 ;
 END
END DIB14
PIN DOB14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3171.980 1710.800 3173.100 1711.920 ;
  LAYER metal4 ;
  RECT 3171.980 1710.800 3173.100 1711.920 ;
  LAYER metal3 ;
  RECT 3171.980 1710.800 3173.100 1711.920 ;
  LAYER metal2 ;
  RECT 3171.980 1710.800 3173.100 1711.920 ;
  LAYER metal1 ;
  RECT 3171.980 1710.800 3173.100 1711.920 ;
 END
END DOB14
PIN DIB13
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2780.140 1710.800 2781.260 1711.920 ;
  LAYER metal4 ;
  RECT 2780.140 1710.800 2781.260 1711.920 ;
  LAYER metal3 ;
  RECT 2780.140 1710.800 2781.260 1711.920 ;
  LAYER metal2 ;
  RECT 2780.140 1710.800 2781.260 1711.920 ;
  LAYER metal1 ;
  RECT 2780.140 1710.800 2781.260 1711.920 ;
 END
END DIB13
PIN DOB13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2767.120 1710.800 2768.240 1711.920 ;
  LAYER metal4 ;
  RECT 2767.120 1710.800 2768.240 1711.920 ;
  LAYER metal3 ;
  RECT 2767.120 1710.800 2768.240 1711.920 ;
  LAYER metal2 ;
  RECT 2767.120 1710.800 2768.240 1711.920 ;
  LAYER metal1 ;
  RECT 2767.120 1710.800 2768.240 1711.920 ;
 END
END DOB13
PIN DIB12
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2753.480 1710.800 2754.600 1711.920 ;
  LAYER metal4 ;
  RECT 2753.480 1710.800 2754.600 1711.920 ;
  LAYER metal3 ;
  RECT 2753.480 1710.800 2754.600 1711.920 ;
  LAYER metal2 ;
  RECT 2753.480 1710.800 2754.600 1711.920 ;
  LAYER metal1 ;
  RECT 2753.480 1710.800 2754.600 1711.920 ;
 END
END DIB12
PIN DOB12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2739.840 1710.800 2740.960 1711.920 ;
  LAYER metal4 ;
  RECT 2739.840 1710.800 2740.960 1711.920 ;
  LAYER metal3 ;
  RECT 2739.840 1710.800 2740.960 1711.920 ;
  LAYER metal2 ;
  RECT 2739.840 1710.800 2740.960 1711.920 ;
  LAYER metal1 ;
  RECT 2739.840 1710.800 2740.960 1711.920 ;
 END
END DOB12
PIN DIB11
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2348.000 1710.800 2349.120 1711.920 ;
  LAYER metal4 ;
  RECT 2348.000 1710.800 2349.120 1711.920 ;
  LAYER metal3 ;
  RECT 2348.000 1710.800 2349.120 1711.920 ;
  LAYER metal2 ;
  RECT 2348.000 1710.800 2349.120 1711.920 ;
  LAYER metal1 ;
  RECT 2348.000 1710.800 2349.120 1711.920 ;
 END
END DIB11
PIN DOB11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2334.360 1710.800 2335.480 1711.920 ;
  LAYER metal4 ;
  RECT 2334.360 1710.800 2335.480 1711.920 ;
  LAYER metal3 ;
  RECT 2334.360 1710.800 2335.480 1711.920 ;
  LAYER metal2 ;
  RECT 2334.360 1710.800 2335.480 1711.920 ;
  LAYER metal1 ;
  RECT 2334.360 1710.800 2335.480 1711.920 ;
 END
END DOB11
PIN DIB10
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2321.340 1710.800 2322.460 1711.920 ;
  LAYER metal4 ;
  RECT 2321.340 1710.800 2322.460 1711.920 ;
  LAYER metal3 ;
  RECT 2321.340 1710.800 2322.460 1711.920 ;
  LAYER metal2 ;
  RECT 2321.340 1710.800 2322.460 1711.920 ;
  LAYER metal1 ;
  RECT 2321.340 1710.800 2322.460 1711.920 ;
 END
END DIB10
PIN DOB10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2307.700 1710.800 2308.820 1711.920 ;
  LAYER metal4 ;
  RECT 2307.700 1710.800 2308.820 1711.920 ;
  LAYER metal3 ;
  RECT 2307.700 1710.800 2308.820 1711.920 ;
  LAYER metal2 ;
  RECT 2307.700 1710.800 2308.820 1711.920 ;
  LAYER metal1 ;
  RECT 2307.700 1710.800 2308.820 1711.920 ;
 END
END DOB10
PIN DIB9
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1915.860 1710.800 1916.980 1711.920 ;
  LAYER metal4 ;
  RECT 1915.860 1710.800 1916.980 1711.920 ;
  LAYER metal3 ;
  RECT 1915.860 1710.800 1916.980 1711.920 ;
  LAYER metal2 ;
  RECT 1915.860 1710.800 1916.980 1711.920 ;
  LAYER metal1 ;
  RECT 1915.860 1710.800 1916.980 1711.920 ;
 END
END DIB9
PIN DOB9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1902.220 1710.800 1903.340 1711.920 ;
  LAYER metal4 ;
  RECT 1902.220 1710.800 1903.340 1711.920 ;
  LAYER metal3 ;
  RECT 1902.220 1710.800 1903.340 1711.920 ;
  LAYER metal2 ;
  RECT 1902.220 1710.800 1903.340 1711.920 ;
  LAYER metal1 ;
  RECT 1902.220 1710.800 1903.340 1711.920 ;
 END
END DOB9
PIN DIB8
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1888.580 1710.800 1889.700 1711.920 ;
  LAYER metal4 ;
  RECT 1888.580 1710.800 1889.700 1711.920 ;
  LAYER metal3 ;
  RECT 1888.580 1710.800 1889.700 1711.920 ;
  LAYER metal2 ;
  RECT 1888.580 1710.800 1889.700 1711.920 ;
  LAYER metal1 ;
  RECT 1888.580 1710.800 1889.700 1711.920 ;
 END
END DIB8
PIN DOB8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1875.560 1710.800 1876.680 1711.920 ;
  LAYER metal4 ;
  RECT 1875.560 1710.800 1876.680 1711.920 ;
  LAYER metal3 ;
  RECT 1875.560 1710.800 1876.680 1711.920 ;
  LAYER metal2 ;
  RECT 1875.560 1710.800 1876.680 1711.920 ;
  LAYER metal1 ;
  RECT 1875.560 1710.800 1876.680 1711.920 ;
 END
END DOB8
PIN OEB
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1848.280 1710.800 1849.400 1711.920 ;
  LAYER metal4 ;
  RECT 1848.280 1710.800 1849.400 1711.920 ;
  LAYER metal3 ;
  RECT 1848.280 1710.800 1849.400 1711.920 ;
  LAYER metal2 ;
  RECT 1848.280 1710.800 1849.400 1711.920 ;
  LAYER metal1 ;
  RECT 1848.280 1710.800 1849.400 1711.920 ;
 END
END OEB
PIN B5
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1843.940 1710.800 1845.060 1711.920 ;
  LAYER metal4 ;
  RECT 1843.940 1710.800 1845.060 1711.920 ;
  LAYER metal3 ;
  RECT 1843.940 1710.800 1845.060 1711.920 ;
  LAYER metal2 ;
  RECT 1843.940 1710.800 1845.060 1711.920 ;
  LAYER metal1 ;
  RECT 1843.940 1710.800 1845.060 1711.920 ;
 END
END B5
PIN B4
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1842.080 1710.800 1843.200 1711.920 ;
  LAYER metal4 ;
  RECT 1842.080 1710.800 1843.200 1711.920 ;
  LAYER metal3 ;
  RECT 1842.080 1710.800 1843.200 1711.920 ;
  LAYER metal2 ;
  RECT 1842.080 1710.800 1843.200 1711.920 ;
  LAYER metal1 ;
  RECT 1842.080 1710.800 1843.200 1711.920 ;
 END
END B4
PIN B3
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1837.120 1710.800 1838.240 1711.920 ;
  LAYER metal4 ;
  RECT 1837.120 1710.800 1838.240 1711.920 ;
  LAYER metal3 ;
  RECT 1837.120 1710.800 1838.240 1711.920 ;
  LAYER metal2 ;
  RECT 1837.120 1710.800 1838.240 1711.920 ;
  LAYER metal1 ;
  RECT 1837.120 1710.800 1838.240 1711.920 ;
 END
END B3
PIN CKB
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1835.260 1710.800 1836.380 1711.920 ;
  LAYER metal4 ;
  RECT 1835.260 1710.800 1836.380 1711.920 ;
  LAYER metal3 ;
  RECT 1835.260 1710.800 1836.380 1711.920 ;
  LAYER metal2 ;
  RECT 1835.260 1710.800 1836.380 1711.920 ;
  LAYER metal1 ;
  RECT 1835.260 1710.800 1836.380 1711.920 ;
 END
END CKB
PIN CSB
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1833.400 1710.800 1834.520 1711.920 ;
  LAYER metal4 ;
  RECT 1833.400 1710.800 1834.520 1711.920 ;
  LAYER metal3 ;
  RECT 1833.400 1710.800 1834.520 1711.920 ;
  LAYER metal2 ;
  RECT 1833.400 1710.800 1834.520 1711.920 ;
  LAYER metal1 ;
  RECT 1833.400 1710.800 1834.520 1711.920 ;
 END
END CSB
PIN WEBN
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1830.300 1710.800 1831.420 1711.920 ;
  LAYER metal4 ;
  RECT 1830.300 1710.800 1831.420 1711.920 ;
  LAYER metal3 ;
  RECT 1830.300 1710.800 1831.420 1711.920 ;
  LAYER metal2 ;
  RECT 1830.300 1710.800 1831.420 1711.920 ;
  LAYER metal1 ;
  RECT 1830.300 1710.800 1831.420 1711.920 ;
 END
END WEBN
PIN B2
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1826.580 1710.800 1827.700 1711.920 ;
  LAYER metal4 ;
  RECT 1826.580 1710.800 1827.700 1711.920 ;
  LAYER metal3 ;
  RECT 1826.580 1710.800 1827.700 1711.920 ;
  LAYER metal2 ;
  RECT 1826.580 1710.800 1827.700 1711.920 ;
  LAYER metal1 ;
  RECT 1826.580 1710.800 1827.700 1711.920 ;
 END
END B2
PIN B1
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1821.620 1710.800 1822.740 1711.920 ;
  LAYER metal4 ;
  RECT 1821.620 1710.800 1822.740 1711.920 ;
  LAYER metal3 ;
  RECT 1821.620 1710.800 1822.740 1711.920 ;
  LAYER metal2 ;
  RECT 1821.620 1710.800 1822.740 1711.920 ;
  LAYER metal1 ;
  RECT 1821.620 1710.800 1822.740 1711.920 ;
 END
END B1
PIN B0
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1819.140 1710.800 1820.260 1711.920 ;
  LAYER metal4 ;
  RECT 1819.140 1710.800 1820.260 1711.920 ;
  LAYER metal3 ;
  RECT 1819.140 1710.800 1820.260 1711.920 ;
  LAYER metal2 ;
  RECT 1819.140 1710.800 1820.260 1711.920 ;
  LAYER metal1 ;
  RECT 1819.140 1710.800 1820.260 1711.920 ;
 END
END B0
PIN B8
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1811.080 1710.800 1812.200 1711.920 ;
  LAYER metal4 ;
  RECT 1811.080 1710.800 1812.200 1711.920 ;
  LAYER metal3 ;
  RECT 1811.080 1710.800 1812.200 1711.920 ;
  LAYER metal2 ;
  RECT 1811.080 1710.800 1812.200 1711.920 ;
  LAYER metal1 ;
  RECT 1811.080 1710.800 1812.200 1711.920 ;
 END
END B8
PIN B7
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1805.500 1710.800 1806.620 1711.920 ;
  LAYER metal4 ;
  RECT 1805.500 1710.800 1806.620 1711.920 ;
  LAYER metal3 ;
  RECT 1805.500 1710.800 1806.620 1711.920 ;
  LAYER metal2 ;
  RECT 1805.500 1710.800 1806.620 1711.920 ;
  LAYER metal1 ;
  RECT 1805.500 1710.800 1806.620 1711.920 ;
 END
END B7
PIN B6
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1799.300 1710.800 1800.420 1711.920 ;
  LAYER metal4 ;
  RECT 1799.300 1710.800 1800.420 1711.920 ;
  LAYER metal3 ;
  RECT 1799.300 1710.800 1800.420 1711.920 ;
  LAYER metal2 ;
  RECT 1799.300 1710.800 1800.420 1711.920 ;
  LAYER metal1 ;
  RECT 1799.300 1710.800 1800.420 1711.920 ;
 END
END B6
PIN B11
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1786.900 1710.800 1788.020 1711.920 ;
  LAYER metal4 ;
  RECT 1786.900 1710.800 1788.020 1711.920 ;
  LAYER metal3 ;
  RECT 1786.900 1710.800 1788.020 1711.920 ;
  LAYER metal2 ;
  RECT 1786.900 1710.800 1788.020 1711.920 ;
  LAYER metal1 ;
  RECT 1786.900 1710.800 1788.020 1711.920 ;
 END
END B11
PIN B10
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1780.700 1710.800 1781.820 1711.920 ;
  LAYER metal4 ;
  RECT 1780.700 1710.800 1781.820 1711.920 ;
  LAYER metal3 ;
  RECT 1780.700 1710.800 1781.820 1711.920 ;
  LAYER metal2 ;
  RECT 1780.700 1710.800 1781.820 1711.920 ;
  LAYER metal1 ;
  RECT 1780.700 1710.800 1781.820 1711.920 ;
 END
END B10
PIN B9
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1775.120 1710.800 1776.240 1711.920 ;
  LAYER metal4 ;
  RECT 1775.120 1710.800 1776.240 1711.920 ;
  LAYER metal3 ;
  RECT 1775.120 1710.800 1776.240 1711.920 ;
  LAYER metal2 ;
  RECT 1775.120 1710.800 1776.240 1711.920 ;
  LAYER metal1 ;
  RECT 1775.120 1710.800 1776.240 1711.920 ;
 END
END B9
PIN B14
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1762.100 1710.800 1763.220 1711.920 ;
  LAYER metal4 ;
  RECT 1762.100 1710.800 1763.220 1711.920 ;
  LAYER metal3 ;
  RECT 1762.100 1710.800 1763.220 1711.920 ;
  LAYER metal2 ;
  RECT 1762.100 1710.800 1763.220 1711.920 ;
  LAYER metal1 ;
  RECT 1762.100 1710.800 1763.220 1711.920 ;
 END
END B14
PIN B13
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1756.520 1710.800 1757.640 1711.920 ;
  LAYER metal4 ;
  RECT 1756.520 1710.800 1757.640 1711.920 ;
  LAYER metal3 ;
  RECT 1756.520 1710.800 1757.640 1711.920 ;
  LAYER metal2 ;
  RECT 1756.520 1710.800 1757.640 1711.920 ;
  LAYER metal1 ;
  RECT 1756.520 1710.800 1757.640 1711.920 ;
 END
END B13
PIN B12
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1750.940 1710.800 1752.060 1711.920 ;
  LAYER metal4 ;
  RECT 1750.940 1710.800 1752.060 1711.920 ;
  LAYER metal3 ;
  RECT 1750.940 1710.800 1752.060 1711.920 ;
  LAYER metal2 ;
  RECT 1750.940 1710.800 1752.060 1711.920 ;
  LAYER metal1 ;
  RECT 1750.940 1710.800 1752.060 1711.920 ;
 END
END B12
PIN DIB7
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1349.800 1710.800 1350.920 1711.920 ;
  LAYER metal4 ;
  RECT 1349.800 1710.800 1350.920 1711.920 ;
  LAYER metal3 ;
  RECT 1349.800 1710.800 1350.920 1711.920 ;
  LAYER metal2 ;
  RECT 1349.800 1710.800 1350.920 1711.920 ;
  LAYER metal1 ;
  RECT 1349.800 1710.800 1350.920 1711.920 ;
 END
END DIB7
PIN DOB7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1336.780 1710.800 1337.900 1711.920 ;
  LAYER metal4 ;
  RECT 1336.780 1710.800 1337.900 1711.920 ;
  LAYER metal3 ;
  RECT 1336.780 1710.800 1337.900 1711.920 ;
  LAYER metal2 ;
  RECT 1336.780 1710.800 1337.900 1711.920 ;
  LAYER metal1 ;
  RECT 1336.780 1710.800 1337.900 1711.920 ;
 END
END DOB7
PIN DIB6
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1323.140 1710.800 1324.260 1711.920 ;
  LAYER metal4 ;
  RECT 1323.140 1710.800 1324.260 1711.920 ;
  LAYER metal3 ;
  RECT 1323.140 1710.800 1324.260 1711.920 ;
  LAYER metal2 ;
  RECT 1323.140 1710.800 1324.260 1711.920 ;
  LAYER metal1 ;
  RECT 1323.140 1710.800 1324.260 1711.920 ;
 END
END DIB6
PIN DOB6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1309.500 1710.800 1310.620 1711.920 ;
  LAYER metal4 ;
  RECT 1309.500 1710.800 1310.620 1711.920 ;
  LAYER metal3 ;
  RECT 1309.500 1710.800 1310.620 1711.920 ;
  LAYER metal2 ;
  RECT 1309.500 1710.800 1310.620 1711.920 ;
  LAYER metal1 ;
  RECT 1309.500 1710.800 1310.620 1711.920 ;
 END
END DOB6
PIN DIB5
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 917.660 1710.800 918.780 1711.920 ;
  LAYER metal4 ;
  RECT 917.660 1710.800 918.780 1711.920 ;
  LAYER metal3 ;
  RECT 917.660 1710.800 918.780 1711.920 ;
  LAYER metal2 ;
  RECT 917.660 1710.800 918.780 1711.920 ;
  LAYER metal1 ;
  RECT 917.660 1710.800 918.780 1711.920 ;
 END
END DIB5
PIN DOB5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 904.020 1710.800 905.140 1711.920 ;
  LAYER metal4 ;
  RECT 904.020 1710.800 905.140 1711.920 ;
  LAYER metal3 ;
  RECT 904.020 1710.800 905.140 1711.920 ;
  LAYER metal2 ;
  RECT 904.020 1710.800 905.140 1711.920 ;
  LAYER metal1 ;
  RECT 904.020 1710.800 905.140 1711.920 ;
 END
END DOB5
PIN DIB4
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 891.000 1710.800 892.120 1711.920 ;
  LAYER metal4 ;
  RECT 891.000 1710.800 892.120 1711.920 ;
  LAYER metal3 ;
  RECT 891.000 1710.800 892.120 1711.920 ;
  LAYER metal2 ;
  RECT 891.000 1710.800 892.120 1711.920 ;
  LAYER metal1 ;
  RECT 891.000 1710.800 892.120 1711.920 ;
 END
END DIB4
PIN DOB4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 877.360 1710.800 878.480 1711.920 ;
  LAYER metal4 ;
  RECT 877.360 1710.800 878.480 1711.920 ;
  LAYER metal3 ;
  RECT 877.360 1710.800 878.480 1711.920 ;
  LAYER metal2 ;
  RECT 877.360 1710.800 878.480 1711.920 ;
  LAYER metal1 ;
  RECT 877.360 1710.800 878.480 1711.920 ;
 END
END DOB4
PIN DIB3
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 485.520 1710.800 486.640 1711.920 ;
  LAYER metal4 ;
  RECT 485.520 1710.800 486.640 1711.920 ;
  LAYER metal3 ;
  RECT 485.520 1710.800 486.640 1711.920 ;
  LAYER metal2 ;
  RECT 485.520 1710.800 486.640 1711.920 ;
  LAYER metal1 ;
  RECT 485.520 1710.800 486.640 1711.920 ;
 END
END DIB3
PIN DOB3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 471.880 1710.800 473.000 1711.920 ;
  LAYER metal4 ;
  RECT 471.880 1710.800 473.000 1711.920 ;
  LAYER metal3 ;
  RECT 471.880 1710.800 473.000 1711.920 ;
  LAYER metal2 ;
  RECT 471.880 1710.800 473.000 1711.920 ;
  LAYER metal1 ;
  RECT 471.880 1710.800 473.000 1711.920 ;
 END
END DOB3
PIN DIB2
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 458.240 1710.800 459.360 1711.920 ;
  LAYER metal4 ;
  RECT 458.240 1710.800 459.360 1711.920 ;
  LAYER metal3 ;
  RECT 458.240 1710.800 459.360 1711.920 ;
  LAYER metal2 ;
  RECT 458.240 1710.800 459.360 1711.920 ;
  LAYER metal1 ;
  RECT 458.240 1710.800 459.360 1711.920 ;
 END
END DIB2
PIN DOB2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 445.220 1710.800 446.340 1711.920 ;
  LAYER metal4 ;
  RECT 445.220 1710.800 446.340 1711.920 ;
  LAYER metal3 ;
  RECT 445.220 1710.800 446.340 1711.920 ;
  LAYER metal2 ;
  RECT 445.220 1710.800 446.340 1711.920 ;
  LAYER metal1 ;
  RECT 445.220 1710.800 446.340 1711.920 ;
 END
END DOB2
PIN DIB1
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 52.760 1710.800 53.880 1711.920 ;
  LAYER metal4 ;
  RECT 52.760 1710.800 53.880 1711.920 ;
  LAYER metal3 ;
  RECT 52.760 1710.800 53.880 1711.920 ;
  LAYER metal2 ;
  RECT 52.760 1710.800 53.880 1711.920 ;
  LAYER metal1 ;
  RECT 52.760 1710.800 53.880 1711.920 ;
 END
END DIB1
PIN DOB1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 39.740 1710.800 40.860 1711.920 ;
  LAYER metal4 ;
  RECT 39.740 1710.800 40.860 1711.920 ;
  LAYER metal3 ;
  RECT 39.740 1710.800 40.860 1711.920 ;
  LAYER metal2 ;
  RECT 39.740 1710.800 40.860 1711.920 ;
  LAYER metal1 ;
  RECT 39.740 1710.800 40.860 1711.920 ;
 END
END DOB1
PIN DIB0
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 26.100 1710.800 27.220 1711.920 ;
  LAYER metal4 ;
  RECT 26.100 1710.800 27.220 1711.920 ;
  LAYER metal3 ;
  RECT 26.100 1710.800 27.220 1711.920 ;
  LAYER metal2 ;
  RECT 26.100 1710.800 27.220 1711.920 ;
  LAYER metal1 ;
  RECT 26.100 1710.800 27.220 1711.920 ;
 END
END DIB0
PIN DOB0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 12.460 1710.800 13.580 1711.920 ;
  LAYER metal4 ;
  RECT 12.460 1710.800 13.580 1711.920 ;
  LAYER metal3 ;
  RECT 12.460 1710.800 13.580 1711.920 ;
  LAYER metal2 ;
  RECT 12.460 1710.800 13.580 1711.920 ;
  LAYER metal1 ;
  RECT 12.460 1710.800 13.580 1711.920 ;
 END
END DOB0
PIN DIA15
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3212.280 0.000 3213.400 1.120 ;
  LAYER metal4 ;
  RECT 3212.280 0.000 3213.400 1.120 ;
  LAYER metal3 ;
  RECT 3212.280 0.000 3213.400 1.120 ;
  LAYER metal2 ;
  RECT 3212.280 0.000 3213.400 1.120 ;
  LAYER metal1 ;
  RECT 3212.280 0.000 3213.400 1.120 ;
 END
END DIA15
PIN DOA15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3199.260 0.000 3200.380 1.120 ;
  LAYER metal4 ;
  RECT 3199.260 0.000 3200.380 1.120 ;
  LAYER metal3 ;
  RECT 3199.260 0.000 3200.380 1.120 ;
  LAYER metal2 ;
  RECT 3199.260 0.000 3200.380 1.120 ;
  LAYER metal1 ;
  RECT 3199.260 0.000 3200.380 1.120 ;
 END
END DOA15
PIN DIA14
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3185.620 0.000 3186.740 1.120 ;
  LAYER metal4 ;
  RECT 3185.620 0.000 3186.740 1.120 ;
  LAYER metal3 ;
  RECT 3185.620 0.000 3186.740 1.120 ;
  LAYER metal2 ;
  RECT 3185.620 0.000 3186.740 1.120 ;
  LAYER metal1 ;
  RECT 3185.620 0.000 3186.740 1.120 ;
 END
END DIA14
PIN DOA14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3171.980 0.000 3173.100 1.120 ;
  LAYER metal4 ;
  RECT 3171.980 0.000 3173.100 1.120 ;
  LAYER metal3 ;
  RECT 3171.980 0.000 3173.100 1.120 ;
  LAYER metal2 ;
  RECT 3171.980 0.000 3173.100 1.120 ;
  LAYER metal1 ;
  RECT 3171.980 0.000 3173.100 1.120 ;
 END
END DOA14
PIN DIA13
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2780.140 0.000 2781.260 1.120 ;
  LAYER metal4 ;
  RECT 2780.140 0.000 2781.260 1.120 ;
  LAYER metal3 ;
  RECT 2780.140 0.000 2781.260 1.120 ;
  LAYER metal2 ;
  RECT 2780.140 0.000 2781.260 1.120 ;
  LAYER metal1 ;
  RECT 2780.140 0.000 2781.260 1.120 ;
 END
END DIA13
PIN DOA13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2767.120 0.000 2768.240 1.120 ;
  LAYER metal4 ;
  RECT 2767.120 0.000 2768.240 1.120 ;
  LAYER metal3 ;
  RECT 2767.120 0.000 2768.240 1.120 ;
  LAYER metal2 ;
  RECT 2767.120 0.000 2768.240 1.120 ;
  LAYER metal1 ;
  RECT 2767.120 0.000 2768.240 1.120 ;
 END
END DOA13
PIN DIA12
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2753.480 0.000 2754.600 1.120 ;
  LAYER metal4 ;
  RECT 2753.480 0.000 2754.600 1.120 ;
  LAYER metal3 ;
  RECT 2753.480 0.000 2754.600 1.120 ;
  LAYER metal2 ;
  RECT 2753.480 0.000 2754.600 1.120 ;
  LAYER metal1 ;
  RECT 2753.480 0.000 2754.600 1.120 ;
 END
END DIA12
PIN DOA12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2739.840 0.000 2740.960 1.120 ;
  LAYER metal4 ;
  RECT 2739.840 0.000 2740.960 1.120 ;
  LAYER metal3 ;
  RECT 2739.840 0.000 2740.960 1.120 ;
  LAYER metal2 ;
  RECT 2739.840 0.000 2740.960 1.120 ;
  LAYER metal1 ;
  RECT 2739.840 0.000 2740.960 1.120 ;
 END
END DOA12
PIN DIA11
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2348.000 0.000 2349.120 1.120 ;
  LAYER metal4 ;
  RECT 2348.000 0.000 2349.120 1.120 ;
  LAYER metal3 ;
  RECT 2348.000 0.000 2349.120 1.120 ;
  LAYER metal2 ;
  RECT 2348.000 0.000 2349.120 1.120 ;
  LAYER metal1 ;
  RECT 2348.000 0.000 2349.120 1.120 ;
 END
END DIA11
PIN DOA11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2334.360 0.000 2335.480 1.120 ;
  LAYER metal4 ;
  RECT 2334.360 0.000 2335.480 1.120 ;
  LAYER metal3 ;
  RECT 2334.360 0.000 2335.480 1.120 ;
  LAYER metal2 ;
  RECT 2334.360 0.000 2335.480 1.120 ;
  LAYER metal1 ;
  RECT 2334.360 0.000 2335.480 1.120 ;
 END
END DOA11
PIN DIA10
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2321.340 0.000 2322.460 1.120 ;
  LAYER metal4 ;
  RECT 2321.340 0.000 2322.460 1.120 ;
  LAYER metal3 ;
  RECT 2321.340 0.000 2322.460 1.120 ;
  LAYER metal2 ;
  RECT 2321.340 0.000 2322.460 1.120 ;
  LAYER metal1 ;
  RECT 2321.340 0.000 2322.460 1.120 ;
 END
END DIA10
PIN DOA10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2307.700 0.000 2308.820 1.120 ;
  LAYER metal4 ;
  RECT 2307.700 0.000 2308.820 1.120 ;
  LAYER metal3 ;
  RECT 2307.700 0.000 2308.820 1.120 ;
  LAYER metal2 ;
  RECT 2307.700 0.000 2308.820 1.120 ;
  LAYER metal1 ;
  RECT 2307.700 0.000 2308.820 1.120 ;
 END
END DOA10
PIN DIA9
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1915.860 0.000 1916.980 1.120 ;
  LAYER metal4 ;
  RECT 1915.860 0.000 1916.980 1.120 ;
  LAYER metal3 ;
  RECT 1915.860 0.000 1916.980 1.120 ;
  LAYER metal2 ;
  RECT 1915.860 0.000 1916.980 1.120 ;
  LAYER metal1 ;
  RECT 1915.860 0.000 1916.980 1.120 ;
 END
END DIA9
PIN DOA9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1902.220 0.000 1903.340 1.120 ;
  LAYER metal4 ;
  RECT 1902.220 0.000 1903.340 1.120 ;
  LAYER metal3 ;
  RECT 1902.220 0.000 1903.340 1.120 ;
  LAYER metal2 ;
  RECT 1902.220 0.000 1903.340 1.120 ;
  LAYER metal1 ;
  RECT 1902.220 0.000 1903.340 1.120 ;
 END
END DOA9
PIN DIA8
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1888.580 0.000 1889.700 1.120 ;
  LAYER metal4 ;
  RECT 1888.580 0.000 1889.700 1.120 ;
  LAYER metal3 ;
  RECT 1888.580 0.000 1889.700 1.120 ;
  LAYER metal2 ;
  RECT 1888.580 0.000 1889.700 1.120 ;
  LAYER metal1 ;
  RECT 1888.580 0.000 1889.700 1.120 ;
 END
END DIA8
PIN DOA8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1875.560 0.000 1876.680 1.120 ;
  LAYER metal4 ;
  RECT 1875.560 0.000 1876.680 1.120 ;
  LAYER metal3 ;
  RECT 1875.560 0.000 1876.680 1.120 ;
  LAYER metal2 ;
  RECT 1875.560 0.000 1876.680 1.120 ;
  LAYER metal1 ;
  RECT 1875.560 0.000 1876.680 1.120 ;
 END
END DOA8
PIN OEA
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1848.280 0.000 1849.400 1.120 ;
  LAYER metal4 ;
  RECT 1848.280 0.000 1849.400 1.120 ;
  LAYER metal3 ;
  RECT 1848.280 0.000 1849.400 1.120 ;
  LAYER metal2 ;
  RECT 1848.280 0.000 1849.400 1.120 ;
  LAYER metal1 ;
  RECT 1848.280 0.000 1849.400 1.120 ;
 END
END OEA
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1843.940 0.000 1845.060 1.120 ;
  LAYER metal4 ;
  RECT 1843.940 0.000 1845.060 1.120 ;
  LAYER metal3 ;
  RECT 1843.940 0.000 1845.060 1.120 ;
  LAYER metal2 ;
  RECT 1843.940 0.000 1845.060 1.120 ;
  LAYER metal1 ;
  RECT 1843.940 0.000 1845.060 1.120 ;
 END
END A5
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1842.080 0.000 1843.200 1.120 ;
  LAYER metal4 ;
  RECT 1842.080 0.000 1843.200 1.120 ;
  LAYER metal3 ;
  RECT 1842.080 0.000 1843.200 1.120 ;
  LAYER metal2 ;
  RECT 1842.080 0.000 1843.200 1.120 ;
  LAYER metal1 ;
  RECT 1842.080 0.000 1843.200 1.120 ;
 END
END A4
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1837.120 0.000 1838.240 1.120 ;
  LAYER metal4 ;
  RECT 1837.120 0.000 1838.240 1.120 ;
  LAYER metal3 ;
  RECT 1837.120 0.000 1838.240 1.120 ;
  LAYER metal2 ;
  RECT 1837.120 0.000 1838.240 1.120 ;
  LAYER metal1 ;
  RECT 1837.120 0.000 1838.240 1.120 ;
 END
END A3
PIN CKA
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1835.260 0.000 1836.380 1.120 ;
  LAYER metal4 ;
  RECT 1835.260 0.000 1836.380 1.120 ;
  LAYER metal3 ;
  RECT 1835.260 0.000 1836.380 1.120 ;
  LAYER metal2 ;
  RECT 1835.260 0.000 1836.380 1.120 ;
  LAYER metal1 ;
  RECT 1835.260 0.000 1836.380 1.120 ;
 END
END CKA
PIN CSA
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1833.400 0.000 1834.520 1.120 ;
  LAYER metal4 ;
  RECT 1833.400 0.000 1834.520 1.120 ;
  LAYER metal3 ;
  RECT 1833.400 0.000 1834.520 1.120 ;
  LAYER metal2 ;
  RECT 1833.400 0.000 1834.520 1.120 ;
  LAYER metal1 ;
  RECT 1833.400 0.000 1834.520 1.120 ;
 END
END CSA
PIN WEAN
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1830.300 0.000 1831.420 1.120 ;
  LAYER metal4 ;
  RECT 1830.300 0.000 1831.420 1.120 ;
  LAYER metal3 ;
  RECT 1830.300 0.000 1831.420 1.120 ;
  LAYER metal2 ;
  RECT 1830.300 0.000 1831.420 1.120 ;
  LAYER metal1 ;
  RECT 1830.300 0.000 1831.420 1.120 ;
 END
END WEAN
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1826.580 0.000 1827.700 1.120 ;
  LAYER metal4 ;
  RECT 1826.580 0.000 1827.700 1.120 ;
  LAYER metal3 ;
  RECT 1826.580 0.000 1827.700 1.120 ;
  LAYER metal2 ;
  RECT 1826.580 0.000 1827.700 1.120 ;
  LAYER metal1 ;
  RECT 1826.580 0.000 1827.700 1.120 ;
 END
END A2
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1821.620 0.000 1822.740 1.120 ;
  LAYER metal4 ;
  RECT 1821.620 0.000 1822.740 1.120 ;
  LAYER metal3 ;
  RECT 1821.620 0.000 1822.740 1.120 ;
  LAYER metal2 ;
  RECT 1821.620 0.000 1822.740 1.120 ;
  LAYER metal1 ;
  RECT 1821.620 0.000 1822.740 1.120 ;
 END
END A1
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1819.140 0.000 1820.260 1.120 ;
  LAYER metal4 ;
  RECT 1819.140 0.000 1820.260 1.120 ;
  LAYER metal3 ;
  RECT 1819.140 0.000 1820.260 1.120 ;
  LAYER metal2 ;
  RECT 1819.140 0.000 1820.260 1.120 ;
  LAYER metal1 ;
  RECT 1819.140 0.000 1820.260 1.120 ;
 END
END A0
PIN A8
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1811.080 0.000 1812.200 1.120 ;
  LAYER metal4 ;
  RECT 1811.080 0.000 1812.200 1.120 ;
  LAYER metal3 ;
  RECT 1811.080 0.000 1812.200 1.120 ;
  LAYER metal2 ;
  RECT 1811.080 0.000 1812.200 1.120 ;
  LAYER metal1 ;
  RECT 1811.080 0.000 1812.200 1.120 ;
 END
END A8
PIN A7
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1805.500 0.000 1806.620 1.120 ;
  LAYER metal4 ;
  RECT 1805.500 0.000 1806.620 1.120 ;
  LAYER metal3 ;
  RECT 1805.500 0.000 1806.620 1.120 ;
  LAYER metal2 ;
  RECT 1805.500 0.000 1806.620 1.120 ;
  LAYER metal1 ;
  RECT 1805.500 0.000 1806.620 1.120 ;
 END
END A7
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1799.300 0.000 1800.420 1.120 ;
  LAYER metal4 ;
  RECT 1799.300 0.000 1800.420 1.120 ;
  LAYER metal3 ;
  RECT 1799.300 0.000 1800.420 1.120 ;
  LAYER metal2 ;
  RECT 1799.300 0.000 1800.420 1.120 ;
  LAYER metal1 ;
  RECT 1799.300 0.000 1800.420 1.120 ;
 END
END A6
PIN A11
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1786.900 0.000 1788.020 1.120 ;
  LAYER metal4 ;
  RECT 1786.900 0.000 1788.020 1.120 ;
  LAYER metal3 ;
  RECT 1786.900 0.000 1788.020 1.120 ;
  LAYER metal2 ;
  RECT 1786.900 0.000 1788.020 1.120 ;
  LAYER metal1 ;
  RECT 1786.900 0.000 1788.020 1.120 ;
 END
END A11
PIN A10
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1780.700 0.000 1781.820 1.120 ;
  LAYER metal4 ;
  RECT 1780.700 0.000 1781.820 1.120 ;
  LAYER metal3 ;
  RECT 1780.700 0.000 1781.820 1.120 ;
  LAYER metal2 ;
  RECT 1780.700 0.000 1781.820 1.120 ;
  LAYER metal1 ;
  RECT 1780.700 0.000 1781.820 1.120 ;
 END
END A10
PIN A9
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1775.120 0.000 1776.240 1.120 ;
  LAYER metal4 ;
  RECT 1775.120 0.000 1776.240 1.120 ;
  LAYER metal3 ;
  RECT 1775.120 0.000 1776.240 1.120 ;
  LAYER metal2 ;
  RECT 1775.120 0.000 1776.240 1.120 ;
  LAYER metal1 ;
  RECT 1775.120 0.000 1776.240 1.120 ;
 END
END A9
PIN A14
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1762.100 0.000 1763.220 1.120 ;
  LAYER metal4 ;
  RECT 1762.100 0.000 1763.220 1.120 ;
  LAYER metal3 ;
  RECT 1762.100 0.000 1763.220 1.120 ;
  LAYER metal2 ;
  RECT 1762.100 0.000 1763.220 1.120 ;
  LAYER metal1 ;
  RECT 1762.100 0.000 1763.220 1.120 ;
 END
END A14
PIN A13
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1756.520 0.000 1757.640 1.120 ;
  LAYER metal4 ;
  RECT 1756.520 0.000 1757.640 1.120 ;
  LAYER metal3 ;
  RECT 1756.520 0.000 1757.640 1.120 ;
  LAYER metal2 ;
  RECT 1756.520 0.000 1757.640 1.120 ;
  LAYER metal1 ;
  RECT 1756.520 0.000 1757.640 1.120 ;
 END
END A13
PIN A12
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1750.940 0.000 1752.060 1.120 ;
  LAYER metal4 ;
  RECT 1750.940 0.000 1752.060 1.120 ;
  LAYER metal3 ;
  RECT 1750.940 0.000 1752.060 1.120 ;
  LAYER metal2 ;
  RECT 1750.940 0.000 1752.060 1.120 ;
  LAYER metal1 ;
  RECT 1750.940 0.000 1752.060 1.120 ;
 END
END A12
PIN DIA7
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1349.800 0.000 1350.920 1.120 ;
  LAYER metal4 ;
  RECT 1349.800 0.000 1350.920 1.120 ;
  LAYER metal3 ;
  RECT 1349.800 0.000 1350.920 1.120 ;
  LAYER metal2 ;
  RECT 1349.800 0.000 1350.920 1.120 ;
  LAYER metal1 ;
  RECT 1349.800 0.000 1350.920 1.120 ;
 END
END DIA7
PIN DOA7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1336.780 0.000 1337.900 1.120 ;
  LAYER metal4 ;
  RECT 1336.780 0.000 1337.900 1.120 ;
  LAYER metal3 ;
  RECT 1336.780 0.000 1337.900 1.120 ;
  LAYER metal2 ;
  RECT 1336.780 0.000 1337.900 1.120 ;
  LAYER metal1 ;
  RECT 1336.780 0.000 1337.900 1.120 ;
 END
END DOA7
PIN DIA6
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1323.140 0.000 1324.260 1.120 ;
  LAYER metal4 ;
  RECT 1323.140 0.000 1324.260 1.120 ;
  LAYER metal3 ;
  RECT 1323.140 0.000 1324.260 1.120 ;
  LAYER metal2 ;
  RECT 1323.140 0.000 1324.260 1.120 ;
  LAYER metal1 ;
  RECT 1323.140 0.000 1324.260 1.120 ;
 END
END DIA6
PIN DOA6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1309.500 0.000 1310.620 1.120 ;
  LAYER metal4 ;
  RECT 1309.500 0.000 1310.620 1.120 ;
  LAYER metal3 ;
  RECT 1309.500 0.000 1310.620 1.120 ;
  LAYER metal2 ;
  RECT 1309.500 0.000 1310.620 1.120 ;
  LAYER metal1 ;
  RECT 1309.500 0.000 1310.620 1.120 ;
 END
END DOA6
PIN DIA5
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 917.660 0.000 918.780 1.120 ;
  LAYER metal4 ;
  RECT 917.660 0.000 918.780 1.120 ;
  LAYER metal3 ;
  RECT 917.660 0.000 918.780 1.120 ;
  LAYER metal2 ;
  RECT 917.660 0.000 918.780 1.120 ;
  LAYER metal1 ;
  RECT 917.660 0.000 918.780 1.120 ;
 END
END DIA5
PIN DOA5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 904.020 0.000 905.140 1.120 ;
  LAYER metal4 ;
  RECT 904.020 0.000 905.140 1.120 ;
  LAYER metal3 ;
  RECT 904.020 0.000 905.140 1.120 ;
  LAYER metal2 ;
  RECT 904.020 0.000 905.140 1.120 ;
  LAYER metal1 ;
  RECT 904.020 0.000 905.140 1.120 ;
 END
END DOA5
PIN DIA4
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 891.000 0.000 892.120 1.120 ;
  LAYER metal4 ;
  RECT 891.000 0.000 892.120 1.120 ;
  LAYER metal3 ;
  RECT 891.000 0.000 892.120 1.120 ;
  LAYER metal2 ;
  RECT 891.000 0.000 892.120 1.120 ;
  LAYER metal1 ;
  RECT 891.000 0.000 892.120 1.120 ;
 END
END DIA4
PIN DOA4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 877.360 0.000 878.480 1.120 ;
  LAYER metal4 ;
  RECT 877.360 0.000 878.480 1.120 ;
  LAYER metal3 ;
  RECT 877.360 0.000 878.480 1.120 ;
  LAYER metal2 ;
  RECT 877.360 0.000 878.480 1.120 ;
  LAYER metal1 ;
  RECT 877.360 0.000 878.480 1.120 ;
 END
END DOA4
PIN DIA3
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 485.520 0.000 486.640 1.120 ;
  LAYER metal4 ;
  RECT 485.520 0.000 486.640 1.120 ;
  LAYER metal3 ;
  RECT 485.520 0.000 486.640 1.120 ;
  LAYER metal2 ;
  RECT 485.520 0.000 486.640 1.120 ;
  LAYER metal1 ;
  RECT 485.520 0.000 486.640 1.120 ;
 END
END DIA3
PIN DOA3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 471.880 0.000 473.000 1.120 ;
  LAYER metal4 ;
  RECT 471.880 0.000 473.000 1.120 ;
  LAYER metal3 ;
  RECT 471.880 0.000 473.000 1.120 ;
  LAYER metal2 ;
  RECT 471.880 0.000 473.000 1.120 ;
  LAYER metal1 ;
  RECT 471.880 0.000 473.000 1.120 ;
 END
END DOA3
PIN DIA2
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 458.240 0.000 459.360 1.120 ;
  LAYER metal4 ;
  RECT 458.240 0.000 459.360 1.120 ;
  LAYER metal3 ;
  RECT 458.240 0.000 459.360 1.120 ;
  LAYER metal2 ;
  RECT 458.240 0.000 459.360 1.120 ;
  LAYER metal1 ;
  RECT 458.240 0.000 459.360 1.120 ;
 END
END DIA2
PIN DOA2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 445.220 0.000 446.340 1.120 ;
  LAYER metal4 ;
  RECT 445.220 0.000 446.340 1.120 ;
  LAYER metal3 ;
  RECT 445.220 0.000 446.340 1.120 ;
  LAYER metal2 ;
  RECT 445.220 0.000 446.340 1.120 ;
  LAYER metal1 ;
  RECT 445.220 0.000 446.340 1.120 ;
 END
END DOA2
PIN DIA1
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER metal4 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER metal3 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER metal2 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER metal1 ;
  RECT 52.760 0.000 53.880 1.120 ;
 END
END DIA1
PIN DOA1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER metal4 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER metal3 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER metal2 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER metal1 ;
  RECT 39.740 0.000 40.860 1.120 ;
 END
END DOA1
PIN DIA0
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER metal4 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER metal3 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER metal2 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER metal1 ;
  RECT 26.100 0.000 27.220 1.120 ;
 END
END DIA0
PIN DOA0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER metal4 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER metal3 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER metal2 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER metal1 ;
  RECT 12.460 0.000 13.580 1.120 ;
 END
END DOA0
OBS
  LAYER metal1 SPACING 0.280 ;
  RECT 0.000 0.140 3613.980 1711.780 ;
  LAYER metal2 SPACING 0.320 ;
  RECT 0.000 0.140 3613.980 1711.780 ;
  LAYER metal3 SPACING 0.320 ;
  RECT 0.000 0.140 3613.980 1711.780 ;
  LAYER metal4 SPACING 0.600 ;
  RECT 0.000 0.140 3613.980 1711.780 ;
  LAYER via ;
  RECT 0.000 0.140 3613.980 1711.780 ;
  LAYER via2 ;
  RECT 0.000 0.140 3613.980 1711.780 ;
  LAYER via3 ;
  RECT 0.000 0.140 3613.980 1711.780 ;
END
END SJMA180_32768X16X1BM8
END LIBRARY



