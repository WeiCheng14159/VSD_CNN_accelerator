`ifndef __EPUDEF__
`define __EPUDEF__

    `define EPU_DATA_BITS 32
    `define EPU_ADDR_BITS 32

`endif